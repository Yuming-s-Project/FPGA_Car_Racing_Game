`timescale 1ns / 1ps
module song1(
input clk,reset,pause,
output reg aud_on, wire pwm);

reg [7:0] duty;
reg [14:0] sample;
reg [13:0] counter;

always@(posedge clk)
begin
if(reset | pause)
    begin
    counter<=0;
    sample<=0;
    aud_on <=0;
    end
else
    begin
    aud_on<=1;
    //8000/100M
    counter <= counter + 1; 
    if(&counter)
    sample <= sample + 1;
    end
end


PWM mypwm(clk,duty,pwm);

//bitmap for 4 seconds of Engine Sound sampled at 8000 samples/seconds, 
//8 bit resolution
//used Audacity to conver the sound clip to 
//unsigned 8 bit raw music, then used 
//Bin2h to convert the file int C header.
//C# code for the bitmap,
/*
int main()
{
    //format
	//15'd0: duty=119; 15'd1: duty=135; ... 15'd7: duty=143;
	//sounddata is an int[] defined in a header created using bin2h

	for (int i = 0; i < 2*16384; i += 8) {
		cout << "15'd" << i     << ": duty=" << (int)sounddata[i] << "; ";
		cout << "15'd" << i + 1 << ": duty=" << (int)sounddata[i + 1] << "; ";
		cout << "15'd" << i + 2 << ": duty=" << (int)sounddata[i + 2] << "; ";
		cout << "15'd" << i + 3 << ": duty=" << (int)sounddata[i + 3] << "; ";
		cout << "15'd" << i + 4 << ": duty=" << (int)sounddata[i + 4] << "; ";
		cout << "15'd" << i + 5 << ": duty=" << (int)sounddata[i + 5] << "; ";
		cout << "15'd" << i + 6 << ": duty=" << (int)sounddata[i + 6] << "; ";
		cout << "15'd" << i + 7 << ": duty=" << (int)sounddata[i + 7] << "; " << endl;
	}
	
    return 0;
}
*/
always@*
case(sample)
15'd0: duty=119; 15'd1: duty=135; 15'd2: duty=131; 15'd3: duty=116; 15'd4: duty=122; 15'd5: duty=135; 15'd6: duty=131; 15'd7: duty=143;
15'd8: duty=149; 15'd9: duty=142; 15'd10: duty=137; 15'd11: duty=127; 15'd12: duty=128; 15'd13: duty=142; 15'd14: duty=152; 15'd15: duty=122;
15'd16: duty=125; 15'd17: duty=145; 15'd18: duty=156; 15'd19: duty=155; 15'd20: duty=156; 15'd21: duty=153; 15'd22: duty=154; 15'd23: duty=156;
15'd24: duty=148; 15'd25: duty=160; 15'd26: duty=151; 15'd27: duty=138; 15'd28: duty=125; 15'd29: duty=124; 15'd30: duty=129; 15'd31: duty=142;
15'd32: duty=145; 15'd33: duty=128; 15'd34: duty=126; 15'd35: duty=132; 15'd36: duty=125; 15'd37: duty=120; 15'd38: duty=119; 15'd39: duty=105;
15'd40: duty=105; 15'd41: duty=114; 15'd42: duty=122; 15'd43: duty=116; 15'd44: duty=98; 15'd45: duty=108; 15'd46: duty=117; 15'd47: duty=113;
15'd48: duty=110; 15'd49: duty=121; 15'd50: duty=120; 15'd51: duty=107; 15'd52: duty=108; 15'd53: duty=115; 15'd54: duty=127; 15'd55: duty=132;
15'd56: duty=140; 15'd57: duty=137; 15'd58: duty=130; 15'd59: duty=133; 15'd60: duty=139; 15'd61: duty=131; 15'd62: duty=134; 15'd63: duty=135;
15'd64: duty=125; 15'd65: duty=135; 15'd66: duty=147; 15'd67: duty=146; 15'd68: duty=133; 15'd69: duty=135; 15'd70: duty=141; 15'd71: duty=154;
15'd72: duty=157; 15'd73: duty=138; 15'd74: duty=130; 15'd75: duty=123; 15'd76: duty=123; 15'd77: duty=147; 15'd78: duty=146; 15'd79: duty=146;
15'd80: duty=144; 15'd81: duty=144; 15'd82: duty=153; 15'd83: duty=160; 15'd84: duty=155; 15'd85: duty=141; 15'd86: duty=151; 15'd87: duty=140;
15'd88: duty=130; 15'd89: duty=135; 15'd90: duty=141; 15'd91: duty=127; 15'd92: duty=121; 15'd93: duty=125; 15'd94: duty=144; 15'd95: duty=143;
15'd96: duty=115; 15'd97: duty=108; 15'd98: duty=102; 15'd99: duty=116; 15'd100: duty=104; 15'd101: duty=102; 15'd102: duty=104; 15'd103: duty=99;
15'd104: duty=107; 15'd105: duty=103; 15'd106: duty=120; 15'd107: duty=132; 15'd108: duty=123; 15'd109: duty=123; 15'd110: duty=126; 15'd111: duty=144;
15'd112: duty=149; 15'd113: duty=133; 15'd114: duty=127; 15'd115: duty=108; 15'd116: duty=111; 15'd117: duty=126; 15'd118: duty=125; 15'd119: duty=141;
15'd120: duty=134; 15'd121: duty=122; 15'd122: duty=135; 15'd123: duty=150; 15'd124: duty=149; 15'd125: duty=140; 15'd126: duty=148; 15'd127: duty=145;
15'd128: duty=154; 15'd129: duty=162; 15'd130: duty=153; 15'd131: duty=144; 15'd132: duty=133; 15'd133: duty=139; 15'd134: duty=142; 15'd135: duty=127;
15'd136: duty=131; 15'd137: duty=159; 15'd138: duty=139; 15'd139: duty=132; 15'd140: duty=153; 15'd141: duty=137; 15'd142: duty=130; 15'd143: duty=127;
15'd144: duty=133; 15'd145: duty=137; 15'd146: duty=137; 15'd147: duty=144; 15'd148: duty=149; 15'd149: duty=135; 15'd150: duty=126; 15'd151: duty=120;
15'd152: duty=117; 15'd153: duty=113; 15'd154: duty=111; 15'd155: duty=110; 15'd156: duty=95; 15'd157: duty=107; 15'd158: duty=99; 15'd159: duty=94;
15'd160: duty=93; 15'd161: duty=91; 15'd162: duty=98; 15'd163: duty=105; 15'd164: duty=118; 15'd165: duty=128; 15'd166: duty=120; 15'd167: duty=106;
15'd168: duty=117; 15'd169: duty=129; 15'd170: duty=144; 15'd171: duty=139; 15'd172: duty=139; 15'd173: duty=145; 15'd174: duty=145; 15'd175: duty=153;
15'd176: duty=148; 15'd177: duty=148; 15'd178: duty=123; 15'd179: duty=121; 15'd180: duty=138; 15'd181: duty=149; 15'd182: duty=144; 15'd183: duty=133;
15'd184: duty=134; 15'd185: duty=141; 15'd186: duty=151; 15'd187: duty=147; 15'd188: duty=169; 15'd189: duty=163; 15'd190: duty=157; 15'd191: duty=148;
15'd192: duty=140; 15'd193: duty=132; 15'd194: duty=137; 15'd195: duty=150; 15'd196: duty=149; 15'd197: duty=146; 15'd198: duty=138; 15'd199: duty=145;
15'd200: duty=148; 15'd201: duty=146; 15'd202: duty=144; 15'd203: duty=141; 15'd204: duty=123; 15'd205: duty=126; 15'd206: duty=137; 15'd207: duty=129;
15'd208: duty=117; 15'd209: duty=114; 15'd210: duty=100; 15'd211: duty=106; 15'd212: duty=116; 15'd213: duty=114; 15'd214: duty=108; 15'd215: duty=117;
15'd216: duty=115; 15'd217: duty=89; 15'd218: duty=99; 15'd219: duty=117; 15'd220: duty=116; 15'd221: duty=108; 15'd222: duty=112; 15'd223: duty=123;
15'd224: duty=129; 15'd225: duty=143; 15'd226: duty=153; 15'd227: duty=133; 15'd228: duty=114; 15'd229: duty=120; 15'd230: duty=131; 15'd231: duty=119;
15'd232: duty=115; 15'd233: duty=125; 15'd234: duty=115; 15'd235: duty=124; 15'd236: duty=131; 15'd237: duty=132; 15'd238: duty=141; 15'd239: duty=138;
15'd240: duty=134; 15'd241: duty=137; 15'd242: duty=144; 15'd243: duty=148; 15'd244: duty=150; 15'd245: duty=154; 15'd246: duty=153; 15'd247: duty=149;
15'd248: duty=150; 15'd249: duty=140; 15'd250: duty=135; 15'd251: duty=137; 15'd252: duty=138; 15'd253: duty=145; 15'd254: duty=134; 15'd255: duty=133;
15'd256: duty=144; 15'd257: duty=146; 15'd258: duty=144; 15'd259: duty=147; 15'd260: duty=145; 15'd261: duty=129; 15'd262: duty=119; 15'd263: duty=124;
15'd264: duty=136; 15'd265: duty=129; 15'd266: duty=126; 15'd267: duty=127; 15'd268: duty=112; 15'd269: duty=110; 15'd270: duty=130; 15'd271: duty=122;
15'd272: duty=106; 15'd273: duty=102; 15'd274: duty=112; 15'd275: duty=116; 15'd276: duty=110; 15'd277: duty=127; 15'd278: duty=127; 15'd279: duty=128;
15'd280: duty=131; 15'd281: duty=131; 15'd282: duty=129; 15'd283: duty=124; 15'd284: duty=116; 15'd285: duty=116; 15'd286: duty=122; 15'd287: duty=123;
15'd288: duty=132; 15'd289: duty=127; 15'd290: duty=116; 15'd291: duty=130; 15'd292: duty=135; 15'd293: duty=128; 15'd294: duty=143; 15'd295: duty=151;
15'd296: duty=143; 15'd297: duty=153; 15'd298: duty=151; 15'd299: duty=145; 15'd300: duty=151; 15'd301: duty=133; 15'd302: duty=129; 15'd303: duty=130;
15'd304: duty=140; 15'd305: duty=153; 15'd306: duty=164; 15'd307: duty=153; 15'd308: duty=146; 15'd309: duty=145; 15'd310: duty=125; 15'd311: duty=129;
15'd312: duty=145; 15'd313: duty=140; 15'd314: duty=136; 15'd315: duty=135; 15'd316: duty=128; 15'd317: duty=124; 15'd318: duty=115; 15'd319: duty=115;
15'd320: duty=113; 15'd321: duty=125; 15'd322: duty=123; 15'd323: duty=113; 15'd324: duty=115; 15'd325: duty=118; 15'd326: duty=120; 15'd327: duty=110;
15'd328: duty=114; 15'd329: duty=134; 15'd330: duty=120; 15'd331: duty=110; 15'd332: duty=124; 15'd333: duty=140; 15'd334: duty=138; 15'd335: duty=127;
15'd336: duty=126; 15'd337: duty=131; 15'd338: duty=118; 15'd339: duty=119; 15'd340: duty=124; 15'd341: duty=116; 15'd342: duty=128; 15'd343: duty=120;
15'd344: duty=124; 15'd345: duty=121; 15'd346: duty=129; 15'd347: duty=145; 15'd348: duty=140; 15'd349: duty=135; 15'd350: duty=142; 15'd351: duty=158;
15'd352: duty=150; 15'd353: duty=142; 15'd354: duty=148; 15'd355: duty=142; 15'd356: duty=145; 15'd357: duty=156; 15'd358: duty=151; 15'd359: duty=144;
15'd360: duty=129; 15'd361: duty=129; 15'd362: duty=129; 15'd363: duty=127; 15'd364: duty=137; 15'd365: duty=143; 15'd366: duty=133; 15'd367: duty=121;
15'd368: duty=135; 15'd369: duty=139; 15'd370: duty=137; 15'd371: duty=141; 15'd372: duty=146; 15'd373: duty=155; 15'd374: duty=153; 15'd375: duty=128;
15'd376: duty=105; 15'd377: duty=111; 15'd378: duty=115; 15'd379: duty=107; 15'd380: duty=117; 15'd381: duty=121; 15'd382: duty=114; 15'd383: duty=112;
15'd384: duty=110; 15'd385: duty=116; 15'd386: duty=124; 15'd387: duty=128; 15'd388: duty=112; 15'd389: duty=109; 15'd390: duty=132; 15'd391: duty=146;
15'd392: duty=130; 15'd393: duty=118; 15'd394: duty=121; 15'd395: duty=131; 15'd396: duty=137; 15'd397: duty=129; 15'd398: duty=128; 15'd399: duty=128;
15'd400: duty=137; 15'd401: duty=128; 15'd402: duty=124; 15'd403: duty=136; 15'd404: duty=133; 15'd405: duty=119; 15'd406: duty=124; 15'd407: duty=140;
15'd408: duty=142; 15'd409: duty=143; 15'd410: duty=128; 15'd411: duty=127; 15'd412: duty=138; 15'd413: duty=136; 15'd414: duty=138; 15'd415: duty=148;
15'd416: duty=146; 15'd417: duty=146; 15'd418: duty=151; 15'd419: duty=142; 15'd420: duty=145; 15'd421: duty=142; 15'd422: duty=149; 15'd423: duty=139;
15'd424: duty=145; 15'd425: duty=143; 15'd426: duty=136; 15'd427: duty=154; 15'd428: duty=124; 15'd429: duty=113; 15'd430: duty=128; 15'd431: duty=131;
15'd432: duty=132; 15'd433: duty=131; 15'd434: duty=119; 15'd435: duty=109; 15'd436: duty=101; 15'd437: duty=118; 15'd438: duty=132; 15'd439: duty=127;
15'd440: duty=114; 15'd441: duty=116; 15'd442: duty=135; 15'd443: duty=126; 15'd444: duty=116; 15'd445: duty=121; 15'd446: duty=137; 15'd447: duty=132;
15'd448: duty=109; 15'd449: duty=126; 15'd450: duty=136; 15'd451: duty=122; 15'd452: duty=108; 15'd453: duty=113; 15'd454: duty=131; 15'd455: duty=139;
15'd456: duty=135; 15'd457: duty=126; 15'd458: duty=134; 15'd459: duty=137; 15'd460: duty=133; 15'd461: duty=135; 15'd462: duty=122; 15'd463: duty=115;
15'd464: duty=134; 15'd465: duty=139; 15'd466: duty=140; 15'd467: duty=137; 15'd468: duty=139; 15'd469: duty=145; 15'd470: duty=144; 15'd471: duty=151;
15'd472: duty=164; 15'd473: duty=148; 15'd474: duty=128; 15'd475: duty=120; 15'd476: duty=117; 15'd477: duty=132; 15'd478: duty=133; 15'd479: duty=127;
15'd480: duty=132; 15'd481: duty=139; 15'd482: duty=137; 15'd483: duty=135; 15'd484: duty=135; 15'd485: duty=152; 15'd486: duty=148; 15'd487: duty=131;
15'd488: duty=123; 15'd489: duty=131; 15'd490: duty=133; 15'd491: duty=131; 15'd492: duty=124; 15'd493: duty=116; 15'd494: duty=112; 15'd495: duty=104;
15'd496: duty=107; 15'd497: duty=110; 15'd498: duty=106; 15'd499: duty=116; 15'd500: duty=121; 15'd501: duty=128; 15'd502: duty=141; 15'd503: duty=142;
15'd504: duty=153; 15'd505: duty=139; 15'd506: duty=128; 15'd507: duty=119; 15'd508: duty=122; 15'd509: duty=131; 15'd510: duty=131; 15'd511: duty=133;
15'd512: duty=133; 15'd513: duty=139; 15'd514: duty=138; 15'd515: duty=142; 15'd516: duty=144; 15'd517: duty=143; 15'd518: duty=133; 15'd519: duty=118;
15'd520: duty=128; 15'd521: duty=130; 15'd522: duty=128; 15'd523: duty=131; 15'd524: duty=147; 15'd525: duty=139; 15'd526: duty=121; 15'd527: duty=125;
15'd528: duty=127; 15'd529: duty=132; 15'd530: duty=142; 15'd531: duty=142; 15'd532: duty=128; 15'd533: duty=128; 15'd534: duty=125; 15'd535: duty=131;
15'd536: duty=125; 15'd537: duty=137; 15'd538: duty=141; 15'd539: duty=129; 15'd540: duty=133; 15'd541: duty=127; 15'd542: duty=124; 15'd543: duty=105;
15'd544: duty=107; 15'd545: duty=111; 15'd546: duty=121; 15'd547: duty=121; 15'd548: duty=123; 15'd549: duty=128; 15'd550: duty=114; 15'd551: duty=122;
15'd552: duty=136; 15'd553: duty=134; 15'd554: duty=128; 15'd555: duty=141; 15'd556: duty=139; 15'd557: duty=140; 15'd558: duty=144; 15'd559: duty=141;
15'd560: duty=139; 15'd561: duty=149; 15'd562: duty=151; 15'd563: duty=127; 15'd564: duty=115; 15'd565: duty=113; 15'd566: duty=118; 15'd567: duty=122;
15'd568: duty=133; 15'd569: duty=144; 15'd570: duty=145; 15'd571: duty=134; 15'd572: duty=131; 15'd573: duty=145; 15'd574: duty=145; 15'd575: duty=144;
15'd576: duty=130; 15'd577: duty=121; 15'd578: duty=142; 15'd579: duty=134; 15'd580: duty=137; 15'd581: duty=136; 15'd582: duty=137; 15'd583: duty=141;
15'd584: duty=133; 15'd585: duty=132; 15'd586: duty=122; 15'd587: duty=124; 15'd588: duty=120; 15'd589: duty=115; 15'd590: duty=125; 15'd591: duty=123;
15'd592: duty=122; 15'd593: duty=141; 15'd594: duty=142; 15'd595: duty=145; 15'd596: duty=149; 15'd597: duty=140; 15'd598: duty=138; 15'd599: duty=139;
15'd600: duty=129; 15'd601: duty=112; 15'd602: duty=112; 15'd603: duty=116; 15'd604: duty=119; 15'd605: duty=115; 15'd606: duty=101; 15'd607: duty=101;
15'd608: duty=106; 15'd609: duty=118; 15'd610: duty=125; 15'd611: duty=133; 15'd612: duty=135; 15'd613: duty=130; 15'd614: duty=132; 15'd615: duty=130;
15'd616: duty=145; 15'd617: duty=154; 15'd618: duty=148; 15'd619: duty=134; 15'd620: duty=128; 15'd621: duty=120; 15'd622: duty=127; 15'd623: duty=134;
15'd624: duty=137; 15'd625: duty=146; 15'd626: duty=133; 15'd627: duty=151; 15'd628: duty=159; 15'd629: duty=156; 15'd630: duty=157; 15'd631: duty=137;
15'd632: duty=128; 15'd633: duty=133; 15'd634: duty=131; 15'd635: duty=128; 15'd636: duty=128; 15'd637: duty=116; 15'd638: duty=122; 15'd639: duty=123;
15'd640: duty=127; 15'd641: duty=136; 15'd642: duty=120; 15'd643: duty=122; 15'd644: duty=128; 15'd645: duty=139; 15'd646: duty=145; 15'd647: duty=135;
15'd648: duty=132; 15'd649: duty=134; 15'd650: duty=125; 15'd651: duty=124; 15'd652: duty=140; 15'd653: duty=141; 15'd654: duty=131; 15'd655: duty=118;
15'd656: duty=119; 15'd657: duty=121; 15'd658: duty=111; 15'd659: duty=94; 15'd660: duty=96; 15'd661: duty=123; 15'd662: duty=127; 15'd663: duty=115;
15'd664: duty=114; 15'd665: duty=115; 15'd666: duty=111; 15'd667: duty=116; 15'd668: duty=135; 15'd669: duty=147; 15'd670: duty=146; 15'd671: duty=128;
15'd672: duty=128; 15'd673: duty=135; 15'd674: duty=131; 15'd675: duty=131; 15'd676: duty=123; 15'd677: duty=124; 15'd678: duty=146; 15'd679: duty=155;
15'd680: duty=148; 15'd681: duty=144; 15'd682: duty=126; 15'd683: duty=130; 15'd684: duty=132; 15'd685: duty=133; 15'd686: duty=142; 15'd687: duty=139;
15'd688: duty=160; 15'd689: duty=170; 15'd690: duty=177; 15'd691: duty=179; 15'd692: duty=173; 15'd693: duty=148; 15'd694: duty=123; 15'd695: duty=139;
15'd696: duty=137; 15'd697: duty=130; 15'd698: duty=126; 15'd699: duty=115; 15'd700: duty=124; 15'd701: duty=125; 15'd702: duty=113; 15'd703: duty=109;
15'd704: duty=106; 15'd705: duty=116; 15'd706: duty=116; 15'd707: duty=119; 15'd708: duty=136; 15'd709: duty=137; 15'd710: duty=145; 15'd711: duty=131;
15'd712: duty=109; 15'd713: duty=102; 15'd714: duty=105; 15'd715: duty=105; 15'd716: duty=97; 15'd717: duty=97; 15'd718: duty=113; 15'd719: duty=118;
15'd720: duty=110; 15'd721: duty=125; 15'd722: duty=142; 15'd723: duty=122; 15'd724: duty=125; 15'd725: duty=148; 15'd726: duty=148; 15'd727: duty=143;
15'd728: duty=141; 15'd729: duty=124; 15'd730: duty=117; 15'd731: duty=132; 15'd732: duty=136; 15'd733: duty=135; 15'd734: duty=137; 15'd735: duty=142;
15'd736: duty=145; 15'd737: duty=141; 15'd738: duty=147; 15'd739: duty=160; 15'd740: duty=151; 15'd741: duty=148; 15'd742: duty=142; 15'd743: duty=145;
15'd744: duty=138; 15'd745: duty=134; 15'd746: duty=145; 15'd747: duty=150; 15'd748: duty=143; 15'd749: duty=132; 15'd750: duty=140; 15'd751: duty=132;
15'd752: duty=137; 15'd753: duty=133; 15'd754: duty=119; 15'd755: duty=132; 15'd756: duty=139; 15'd757: duty=140; 15'd758: duty=133; 15'd759: duty=128;
15'd760: duty=125; 15'd761: duty=128; 15'd762: duty=107; 15'd763: duty=89; 15'd764: duty=104; 15'd765: duty=106; 15'd766: duty=121; 15'd767: duty=121;
15'd768: duty=107; 15'd769: duty=107; 15'd770: duty=107; 15'd771: duty=93; 15'd772: duty=98; 15'd773: duty=123; 15'd774: duty=127; 15'd775: duty=121;
15'd776: duty=140; 15'd777: duty=142; 15'd778: duty=140; 15'd779: duty=148; 15'd780: duty=134; 15'd781: duty=127; 15'd782: duty=140; 15'd783: duty=127;
15'd784: duty=118; 15'd785: duty=127; 15'd786: duty=131; 15'd787: duty=140; 15'd788: duty=118; 15'd789: duty=120; 15'd790: duty=145; 15'd791: duty=150;
15'd792: duty=146; 15'd793: duty=148; 15'd794: duty=154; 15'd795: duty=162; 15'd796: duty=167; 15'd797: duty=151; 15'd798: duty=131; 15'd799: duty=130;
15'd800: duty=142; 15'd801: duty=168; 15'd802: duty=163; 15'd803: duty=137; 15'd804: duty=143; 15'd805: duty=139; 15'd806: duty=128; 15'd807: duty=141;
15'd808: duty=142; 15'd809: duty=137; 15'd810: duty=140; 15'd811: duty=145; 15'd812: duty=136; 15'd813: duty=128; 15'd814: duty=113; 15'd815: duty=107;
15'd816: duty=121; 15'd817: duty=124; 15'd818: duty=136; 15'd819: duty=131; 15'd820: duty=115; 15'd821: duty=98; 15'd822: duty=92; 15'd823: duty=87;
15'd824: duty=93; 15'd825: duty=116; 15'd826: duty=128; 15'd827: duty=118; 15'd828: duty=107; 15'd829: duty=110; 15'd830: duty=115; 15'd831: duty=126;
15'd832: duty=128; 15'd833: duty=123; 15'd834: duty=113; 15'd835: duty=134; 15'd836: duty=145; 15'd837: duty=128; 15'd838: duty=121; 15'd839: duty=124;
15'd840: duty=127; 15'd841: duty=129; 15'd842: duty=148; 15'd843: duty=154; 15'd844: duty=145; 15'd845: duty=128; 15'd846: duty=128; 15'd847: duty=130;
15'd848: duty=141; 15'd849: duty=156; 15'd850: duty=167; 15'd851: duty=162; 15'd852: duty=168; 15'd853: duty=173; 15'd854: duty=148; 15'd855: duty=134;
15'd856: duty=128; 15'd857: duty=127; 15'd858: duty=119; 15'd859: duty=131; 15'd860: duty=136; 15'd861: duty=126; 15'd862: duty=131; 15'd863: duty=140;
15'd864: duty=133; 15'd865: duty=134; 15'd866: duty=134; 15'd867: duty=136; 15'd868: duty=134; 15'd869: duty=113; 15'd870: duty=119; 15'd871: duty=125;
15'd872: duty=116; 15'd873: duty=110; 15'd874: duty=112; 15'd875: duty=127; 15'd876: duty=121; 15'd877: duty=115; 15'd878: duty=119; 15'd879: duty=128;
15'd880: duty=127; 15'd881: duty=99; 15'd882: duty=84; 15'd883: duty=110; 15'd884: duty=124; 15'd885: duty=109; 15'd886: duty=113; 15'd887: duty=114;
15'd888: duty=140; 15'd889: duty=153; 15'd890: duty=148; 15'd891: duty=136; 15'd892: duty=128; 15'd893: duty=134; 15'd894: duty=123; 15'd895: duty=132;
15'd896: duty=137; 15'd897: duty=132; 15'd898: duty=123; 15'd899: duty=119; 15'd900: duty=133; 15'd901: duty=155; 15'd902: duty=158; 15'd903: duty=152;
15'd904: duty=149; 15'd905: duty=141; 15'd906: duty=149; 15'd907: duty=141; 15'd908: duty=130; 15'd909: duty=135; 15'd910: duty=136; 15'd911: duty=143;
15'd912: duty=162; 15'd913: duty=169; 15'd914: duty=161; 15'd915: duty=143; 15'd916: duty=135; 15'd917: duty=143; 15'd918: duty=159; 15'd919: duty=164;
15'd920: duty=141; 15'd921: duty=129; 15'd922: duty=119; 15'd923: duty=122; 15'd924: duty=135; 15'd925: duty=143; 15'd926: duty=141; 15'd927: duty=120;
15'd928: duty=121; 15'd929: duty=108; 15'd930: duty=106; 15'd931: duty=109; 15'd932: duty=105; 15'd933: duty=121; 15'd934: duty=124; 15'd935: duty=126;
15'd936: duty=101; 15'd937: duty=100; 15'd938: duty=109; 15'd939: duty=95; 15'd940: duty=89; 15'd941: duty=108; 15'd942: duty=120; 15'd943: duty=114;
15'd944: duty=112; 15'd945: duty=119; 15'd946: duty=122; 15'd947: duty=124; 15'd948: duty=121; 15'd949: duty=115; 15'd950: duty=118; 15'd951: duty=118;
15'd952: duty=126; 15'd953: duty=140; 15'd954: duty=153; 15'd955: duty=148; 15'd956: duty=148; 15'd957: duty=151; 15'd958: duty=154; 15'd959: duty=139;
15'd960: duty=145; 15'd961: duty=147; 15'd962: duty=153; 15'd963: duty=143; 15'd964: duty=134; 15'd965: duty=142; 15'd966: duty=151; 15'd967: duty=151;
15'd968: duty=140; 15'd969: duty=162; 15'd970: duty=151; 15'd971: duty=142; 15'd972: duty=145; 15'd973: duty=150; 15'd974: duty=127; 15'd975: duty=114;
15'd976: duty=110; 15'd977: duty=117; 15'd978: duty=135; 15'd979: duty=156; 15'd980: duty=137; 15'd981: duty=126; 15'd982: duty=122; 15'd983: duty=140;
15'd984: duty=147; 15'd985: duty=123; 15'd986: duty=134; 15'd987: duty=106; 15'd988: duty=119; 15'd989: duty=145; 15'd990: duty=157; 15'd991: duty=131;
15'd992: duty=99; 15'd993: duty=110; 15'd994: duty=104; 15'd995: duty=98; 15'd996: duty=124; 15'd997: duty=124; 15'd998: duty=125; 15'd999: duty=127;
15'd1000: duty=124; 15'd1001: duty=123; 15'd1002: duty=116; 15'd1003: duty=123; 15'd1004: duty=105; 15'd1005: duty=106; 15'd1006: duty=132; 15'd1007: duty=139;
15'd1008: duty=137; 15'd1009: duty=115; 15'd1010: duty=128; 15'd1011: duty=156; 15'd1012: duty=137; 15'd1013: duty=135; 15'd1014: duty=152; 15'd1015: duty=159;
15'd1016: duty=170; 15'd1017: duty=162; 15'd1018: duty=143; 15'd1019: duty=147; 15'd1020: duty=138; 15'd1021: duty=132; 15'd1022: duty=146; 15'd1023: duty=155;
15'd1024: duty=141; 15'd1025: duty=132; 15'd1026: duty=143; 15'd1027: duty=141; 15'd1028: duty=130; 15'd1029: duty=135; 15'd1030: duty=136; 15'd1031: duty=151;
15'd1032: duty=150; 15'd1033: duty=149; 15'd1034: duty=138; 15'd1035: duty=111; 15'd1036: duty=117; 15'd1037: duty=135; 15'd1038: duty=143; 15'd1039: duty=136;
15'd1040: duty=126; 15'd1041: duty=125; 15'd1042: duty=129; 15'd1043: duty=129; 15'd1044: duty=129; 15'd1045: duty=113; 15'd1046: duty=94; 15'd1047: duty=106;
15'd1048: duty=103; 15'd1049: duty=104; 15'd1050: duty=105; 15'd1051: duty=95; 15'd1052: duty=110; 15'd1053: duty=114; 15'd1054: duty=126; 15'd1055: duty=121;
15'd1056: duty=106; 15'd1057: duty=98; 15'd1058: duty=105; 15'd1059: duty=111; 15'd1060: duty=126; 15'd1061: duty=120; 15'd1062: duty=108; 15'd1063: duty=114;
15'd1064: duty=128; 15'd1065: duty=127; 15'd1066: duty=119; 15'd1067: duty=136; 15'd1068: duty=131; 15'd1069: duty=144; 15'd1070: duty=151; 15'd1071: duty=145;
15'd1072: duty=146; 15'd1073: duty=151; 15'd1074: duty=146; 15'd1075: duty=147; 15'd1076: duty=143; 15'd1077: duty=144; 15'd1078: duty=148; 15'd1079: duty=141;
15'd1080: duty=153; 15'd1081: duty=165; 15'd1082: duty=149; 15'd1083: duty=156; 15'd1084: duty=157; 15'd1085: duty=139; 15'd1086: duty=117; 15'd1087: duty=121;
15'd1088: duty=137; 15'd1089: duty=124; 15'd1090: duty=137; 15'd1091: duty=128; 15'd1092: duty=138; 15'd1093: duty=153; 15'd1094: duty=135; 15'd1095: duty=136;
15'd1096: duty=137; 15'd1097: duty=128; 15'd1098: duty=124; 15'd1099: duty=124; 15'd1100: duty=135; 15'd1101: duty=133; 15'd1102: duty=120; 15'd1103: duty=127;
15'd1104: duty=133; 15'd1105: duty=123; 15'd1106: duty=118; 15'd1107: duty=115; 15'd1108: duty=113; 15'd1109: duty=103; 15'd1110: duty=120; 15'd1111: duty=134;
15'd1112: duty=119; 15'd1113: duty=121; 15'd1114: duty=127; 15'd1115: duty=115; 15'd1116: duty=113; 15'd1117: duty=116; 15'd1118: duty=122; 15'd1119: duty=128;
15'd1120: duty=114; 15'd1121: duty=128; 15'd1122: duty=127; 15'd1123: duty=119; 15'd1124: duty=133; 15'd1125: duty=134; 15'd1126: duty=134; 15'd1127: duty=146;
15'd1128: duty=140; 15'd1129: duty=148; 15'd1130: duty=147; 15'd1131: duty=139; 15'd1132: duty=157; 15'd1133: duty=163; 15'd1134: duty=160; 15'd1135: duty=146;
15'd1136: duty=136; 15'd1137: duty=134; 15'd1138: duty=134; 15'd1139: duty=139; 15'd1140: duty=134; 15'd1141: duty=144; 15'd1142: duty=130; 15'd1143: duty=126;
15'd1144: duty=141; 15'd1145: duty=132; 15'd1146: duty=139; 15'd1147: duty=145; 15'd1148: duty=139; 15'd1149: duty=134; 15'd1150: duty=138; 15'd1151: duty=125;
15'd1152: duty=121; 15'd1153: duty=120; 15'd1154: duty=115; 15'd1155: duty=107; 15'd1156: duty=112; 15'd1157: duty=99; 15'd1158: duty=86; 15'd1159: duty=98;
15'd1160: duty=117; 15'd1161: duty=128; 15'd1162: duty=116; 15'd1163: duty=117; 15'd1164: duty=128; 15'd1165: duty=138; 15'd1166: duty=136; 15'd1167: duty=134;
15'd1168: duty=121; 15'd1169: duty=117; 15'd1170: duty=115; 15'd1171: duty=109; 15'd1172: duty=118; 15'd1173: duty=119; 15'd1174: duty=121; 15'd1175: duty=128;
15'd1176: duty=131; 15'd1177: duty=134; 15'd1178: duty=132; 15'd1179: duty=132; 15'd1180: duty=130; 15'd1181: duty=145; 15'd1182: duty=154; 15'd1183: duty=151;
15'd1184: duty=158; 15'd1185: duty=142; 15'd1186: duty=133; 15'd1187: duty=131; 15'd1188: duty=137; 15'd1189: duty=148; 15'd1190: duty=146; 15'd1191: duty=148;
15'd1192: duty=149; 15'd1193: duty=154; 15'd1194: duty=143; 15'd1195: duty=121; 15'd1196: duty=128; 15'd1197: duty=153; 15'd1198: duty=148; 15'd1199: duty=124;
15'd1200: duty=122; 15'd1201: duty=130; 15'd1202: duty=137; 15'd1203: duty=115; 15'd1204: duty=108; 15'd1205: duty=131; 15'd1206: duty=135; 15'd1207: duty=135;
15'd1208: duty=129; 15'd1209: duty=137; 15'd1210: duty=145; 15'd1211: duty=126; 15'd1212: duty=121; 15'd1213: duty=116; 15'd1214: duty=113; 15'd1215: duty=121;
15'd1216: duty=118; 15'd1217: duty=122; 15'd1218: duty=141; 15'd1219: duty=136; 15'd1220: duty=126; 15'd1221: duty=134; 15'd1222: duty=143; 15'd1223: duty=148;
15'd1224: duty=144; 15'd1225: duty=134; 15'd1226: duty=117; 15'd1227: duty=113; 15'd1228: duty=109; 15'd1229: duty=111; 15'd1230: duty=124; 15'd1231: duty=115;
15'd1232: duty=125; 15'd1233: duty=124; 15'd1234: duty=120; 15'd1235: duty=124; 15'd1236: duty=130; 15'd1237: duty=140; 15'd1238: duty=142; 15'd1239: duty=134;
15'd1240: duty=129; 15'd1241: duty=148; 15'd1242: duty=162; 15'd1243: duty=148; 15'd1244: duty=140; 15'd1245: duty=134; 15'd1246: duty=132; 15'd1247: duty=136;
15'd1248: duty=131; 15'd1249: duty=133; 15'd1250: duty=140; 15'd1251: duty=139; 15'd1252: duty=123; 15'd1253: duty=128; 15'd1254: duty=128; 15'd1255: duty=136;
15'd1256: duty=132; 15'd1257: duty=124; 15'd1258: duty=132; 15'd1259: duty=127; 15'd1260: duty=135; 15'd1261: duty=144; 15'd1262: duty=136; 15'd1263: duty=135;
15'd1264: duty=135; 15'd1265: duty=123; 15'd1266: duty=117; 15'd1267: duty=121; 15'd1268: duty=117; 15'd1269: duty=112; 15'd1270: duty=125; 15'd1271: duty=118;
15'd1272: duty=125; 15'd1273: duty=138; 15'd1274: duty=128; 15'd1275: duty=127; 15'd1276: duty=130; 15'd1277: duty=136; 15'd1278: duty=143; 15'd1279: duty=136;
15'd1280: duty=121; 15'd1281: duty=127; 15'd1282: duty=124; 15'd1283: duty=107; 15'd1284: duty=117; 15'd1285: duty=137; 15'd1286: duty=138; 15'd1287: duty=140;
15'd1288: duty=141; 15'd1289: duty=133; 15'd1290: duty=144; 15'd1291: duty=137; 15'd1292: duty=126; 15'd1293: duty=125; 15'd1294: duty=130; 15'd1295: duty=127;
15'd1296: duty=131; 15'd1297: duty=126; 15'd1298: duty=134; 15'd1299: duty=154; 15'd1300: duty=159; 15'd1301: duty=162; 15'd1302: duty=147; 15'd1303: duty=144;
15'd1304: duty=138; 15'd1305: duty=149; 15'd1306: duty=140; 15'd1307: duty=128; 15'd1308: duty=137; 15'd1309: duty=127; 15'd1310: duty=117; 15'd1311: duty=108;
15'd1312: duty=96; 15'd1313: duty=107; 15'd1314: duty=110; 15'd1315: duty=106; 15'd1316: duty=116; 15'd1317: duty=133; 15'd1318: duty=128; 15'd1319: duty=126;
15'd1320: duty=140; 15'd1321: duty=129; 15'd1322: duty=132; 15'd1323: duty=115; 15'd1324: duty=112; 15'd1325: duty=121; 15'd1326: duty=108; 15'd1327: duty=120;
15'd1328: duty=134; 15'd1329: duty=136; 15'd1330: duty=137; 15'd1331: duty=144; 15'd1332: duty=133; 15'd1333: duty=132; 15'd1334: duty=145; 15'd1335: duty=117;
15'd1336: duty=96; 15'd1337: duty=95; 15'd1338: duty=105; 15'd1339: duty=114; 15'd1340: duty=126; 15'd1341: duty=153; 15'd1342: duty=152; 15'd1343: duty=145;
15'd1344: duty=139; 15'd1345: duty=145; 15'd1346: duty=154; 15'd1347: duty=154; 15'd1348: duty=146; 15'd1349: duty=133; 15'd1350: duty=136; 15'd1351: duty=141;
15'd1352: duty=150; 15'd1353: duty=146; 15'd1354: duty=137; 15'd1355: duty=129; 15'd1356: duty=138; 15'd1357: duty=154; 15'd1358: duty=160; 15'd1359: duty=146;
15'd1360: duty=144; 15'd1361: duty=138; 15'd1362: duty=118; 15'd1363: duty=110; 15'd1364: duty=123; 15'd1365: duty=143; 15'd1366: duty=152; 15'd1367: duty=128;
15'd1368: duty=119; 15'd1369: duty=139; 15'd1370: duty=126; 15'd1371: duty=127; 15'd1372: duty=124; 15'd1373: duty=124; 15'd1374: duty=131; 15'd1375: duty=124;
15'd1376: duty=118; 15'd1377: duty=108; 15'd1378: duty=105; 15'd1379: duty=101; 15'd1380: duty=99; 15'd1381: duty=122; 15'd1382: duty=137; 15'd1383: duty=133;
15'd1384: duty=129; 15'd1385: duty=132; 15'd1386: duty=124; 15'd1387: duty=128; 15'd1388: duty=129; 15'd1389: duty=138; 15'd1390: duty=133; 15'd1391: duty=124;
15'd1392: duty=113; 15'd1393: duty=120; 15'd1394: duty=125; 15'd1395: duty=119; 15'd1396: duty=126; 15'd1397: duty=133; 15'd1398: duty=146; 15'd1399: duty=142;
15'd1400: duty=146; 15'd1401: duty=152; 15'd1402: duty=154; 15'd1403: duty=144; 15'd1404: duty=155; 15'd1405: duty=153; 15'd1406: duty=149; 15'd1407: duty=145;
15'd1408: duty=131; 15'd1409: duty=121; 15'd1410: duty=131; 15'd1411: duty=134; 15'd1412: duty=110; 15'd1413: duty=100; 15'd1414: duty=117; 15'd1415: duty=126;
15'd1416: duty=113; 15'd1417: duty=116; 15'd1418: duty=127; 15'd1419: duty=127; 15'd1420: duty=110; 15'd1421: duty=104; 15'd1422: duty=135; 15'd1423: duty=149;
15'd1424: duty=140; 15'd1425: duty=139; 15'd1426: duty=122; 15'd1427: duty=126; 15'd1428: duty=136; 15'd1429: duty=129; 15'd1430: duty=130; 15'd1431: duty=114;
15'd1432: duty=110; 15'd1433: duty=105; 15'd1434: duty=99; 15'd1435: duty=109; 15'd1436: duty=107; 15'd1437: duty=121; 15'd1438: duty=123; 15'd1439: duty=145;
15'd1440: duty=167; 15'd1441: duty=170; 15'd1442: duty=162; 15'd1443: duty=154; 15'd1444: duty=147; 15'd1445: duty=128; 15'd1446: duty=137; 15'd1447: duty=127;
15'd1448: duty=126; 15'd1449: duty=138; 15'd1450: duty=126; 15'd1451: duty=129; 15'd1452: duty=135; 15'd1453: duty=150; 15'd1454: duty=154; 15'd1455: duty=148;
15'd1456: duty=156; 15'd1457: duty=153; 15'd1458: duty=140; 15'd1459: duty=128; 15'd1460: duty=128; 15'd1461: duty=141; 15'd1462: duty=160; 15'd1463: duty=159;
15'd1464: duty=164; 15'd1465: duty=156; 15'd1466: duty=154; 15'd1467: duty=142; 15'd1468: duty=106; 15'd1469: duty=109; 15'd1470: duty=109; 15'd1471: duty=104;
15'd1472: duty=124; 15'd1473: duty=117; 15'd1474: duty=104; 15'd1475: duty=99; 15'd1476: duty=119; 15'd1477: duty=131; 15'd1478: duty=111; 15'd1479: duty=104;
15'd1480: duty=113; 15'd1481: duty=124; 15'd1482: duty=129; 15'd1483: duty=130; 15'd1484: duty=124; 15'd1485: duty=115; 15'd1486: duty=96; 15'd1487: duty=110;
15'd1488: duty=104; 15'd1489: duty=104; 15'd1490: duty=111; 15'd1491: duty=113; 15'd1492: duty=111; 15'd1493: duty=126; 15'd1494: duty=145; 15'd1495: duty=146;
15'd1496: duty=146; 15'd1497: duty=136; 15'd1498: duty=128; 15'd1499: duty=121; 15'd1500: duty=137; 15'd1501: duty=143; 15'd1502: duty=132; 15'd1503: duty=138;
15'd1504: duty=157; 15'd1505: duty=150; 15'd1506: duty=139; 15'd1507: duty=134; 15'd1508: duty=142; 15'd1509: duty=143; 15'd1510: duty=145; 15'd1511: duty=136;
15'd1512: duty=143; 15'd1513: duty=141; 15'd1514: duty=151; 15'd1515: duty=165; 15'd1516: duty=151; 15'd1517: duty=152; 15'd1518: duty=155; 15'd1519: duty=148;
15'd1520: duty=149; 15'd1521: duty=158; 15'd1522: duty=133; 15'd1523: duty=116; 15'd1524: duty=118; 15'd1525: duty=127; 15'd1526: duty=121; 15'd1527: duty=134;
15'd1528: duty=113; 15'd1529: duty=115; 15'd1530: duty=113; 15'd1531: duty=115; 15'd1532: duty=138; 15'd1533: duty=120; 15'd1534: duty=129; 15'd1535: duty=112;
15'd1536: duty=87; 15'd1537: duty=96; 15'd1538: duty=111; 15'd1539: duty=98; 15'd1540: duty=103; 15'd1541: duty=115; 15'd1542: duty=124; 15'd1543: duty=136;
15'd1544: duty=142; 15'd1545: duty=128; 15'd1546: duty=131; 15'd1547: duty=138; 15'd1548: duty=120; 15'd1549: duty=117; 15'd1550: duty=137; 15'd1551: duty=147;
15'd1552: duty=142; 15'd1553: duty=135; 15'd1554: duty=140; 15'd1555: duty=127; 15'd1556: duty=104; 15'd1557: duty=111; 15'd1558: duty=138; 15'd1559: duty=138;
15'd1560: duty=131; 15'd1561: duty=144; 15'd1562: duty=152; 15'd1563: duty=141; 15'd1564: duty=132; 15'd1565: duty=135; 15'd1566: duty=144; 15'd1567: duty=153;
15'd1568: duty=156; 15'd1569: duty=161; 15'd1570: duty=146; 15'd1571: duty=153; 15'd1572: duty=140; 15'd1573: duty=138; 15'd1574: duty=152; 15'd1575: duty=135;
15'd1576: duty=123; 15'd1577: duty=133; 15'd1578: duty=130; 15'd1579: duty=138; 15'd1580: duty=131; 15'd1581: duty=128; 15'd1582: duty=123; 15'd1583: duty=115;
15'd1584: duty=134; 15'd1585: duty=121; 15'd1586: duty=105; 15'd1587: duty=92; 15'd1588: duty=118; 15'd1589: duty=130; 15'd1590: duty=127; 15'd1591: duty=123;
15'd1592: duty=119; 15'd1593: duty=115; 15'd1594: duty=122; 15'd1595: duty=123; 15'd1596: duty=118; 15'd1597: duty=124; 15'd1598: duty=116; 15'd1599: duty=96;
15'd1600: duty=104; 15'd1601: duty=126; 15'd1602: duty=119; 15'd1603: duty=108; 15'd1604: duty=116; 15'd1605: duty=142; 15'd1606: duty=144; 15'd1607: duty=140;
15'd1608: duty=141; 15'd1609: duty=134; 15'd1610: duty=131; 15'd1611: duty=137; 15'd1612: duty=132; 15'd1613: duty=133; 15'd1614: duty=145; 15'd1615: duty=138;
15'd1616: duty=157; 15'd1617: duty=164; 15'd1618: duty=159; 15'd1619: duty=170; 15'd1620: duty=163; 15'd1621: duty=155; 15'd1622: duty=140; 15'd1623: duty=144;
15'd1624: duty=149; 15'd1625: duty=154; 15'd1626: duty=149; 15'd1627: duty=143; 15'd1628: duty=139; 15'd1629: duty=128; 15'd1630: duty=123; 15'd1631: duty=112;
15'd1632: duty=140; 15'd1633: duty=139; 15'd1634: duty=145; 15'd1635: duty=163; 15'd1636: duty=149; 15'd1637: duty=167; 15'd1638: duty=134; 15'd1639: duty=110;
15'd1640: duty=105; 15'd1641: duty=92; 15'd1642: duty=99; 15'd1643: duty=102; 15'd1644: duty=113; 15'd1645: duty=101; 15'd1646: duty=64; 15'd1647: duty=93;
15'd1648: duty=124; 15'd1649: duty=101; 15'd1650: duty=112; 15'd1651: duty=114; 15'd1652: duty=106; 15'd1653: duty=118; 15'd1654: duty=126; 15'd1655: duty=127;
15'd1656: duty=111; 15'd1657: duty=127; 15'd1658: duty=136; 15'd1659: duty=127; 15'd1660: duty=144; 15'd1661: duty=133; 15'd1662: duty=134; 15'd1663: duty=151;
15'd1664: duty=145; 15'd1665: duty=141; 15'd1666: duty=128; 15'd1667: duty=112; 15'd1668: duty=114; 15'd1669: duty=130; 15'd1670: duty=134; 15'd1671: duty=143;
15'd1672: duty=158; 15'd1673: duty=145; 15'd1674: duty=154; 15'd1675: duty=166; 15'd1676: duty=152; 15'd1677: duty=152; 15'd1678: duty=153; 15'd1679: duty=152;
15'd1680: duty=151; 15'd1681: duty=152; 15'd1682: duty=159; 15'd1683: duty=157; 15'd1684: duty=141; 15'd1685: duty=136; 15'd1686: duty=132; 15'd1687: duty=122;
15'd1688: duty=125; 15'd1689: duty=143; 15'd1690: duty=135; 15'd1691: duty=151; 15'd1692: duty=151; 15'd1693: duty=128; 15'd1694: duty=121; 15'd1695: duty=116;
15'd1696: duty=129; 15'd1697: duty=111; 15'd1698: duty=117; 15'd1699: duty=122; 15'd1700: duty=121; 15'd1701: duty=130; 15'd1702: duty=114; 15'd1703: duty=110;
15'd1704: duty=95; 15'd1705: duty=71; 15'd1706: duty=89; 15'd1707: duty=91; 15'd1708: duty=81; 15'd1709: duty=92; 15'd1710: duty=103; 15'd1711: duty=120;
15'd1712: duty=115; 15'd1713: duty=125; 15'd1714: duty=124; 15'd1715: duty=120; 15'd1716: duty=148; 15'd1717: duty=144; 15'd1718: duty=138; 15'd1719: duty=120;
15'd1720: duty=118; 15'd1721: duty=137; 15'd1722: duty=138; 15'd1723: duty=129; 15'd1724: duty=136; 15'd1725: duty=129; 15'd1726: duty=131; 15'd1727: duty=149;
15'd1728: duty=151; 15'd1729: duty=161; 15'd1730: duty=161; 15'd1731: duty=160; 15'd1732: duty=153; 15'd1733: duty=174; 15'd1734: duty=172; 15'd1735: duty=172;
15'd1736: duty=162; 15'd1737: duty=143; 15'd1738: duty=152; 15'd1739: duty=152; 15'd1740: duty=157; 15'd1741: duty=138; 15'd1742: duty=142; 15'd1743: duty=154;
15'd1744: duty=130; 15'd1745: duty=131; 15'd1746: duty=139; 15'd1747: duty=143; 15'd1748: duty=139; 15'd1749: duty=119; 15'd1750: duty=115; 15'd1751: duty=107;
15'd1752: duty=101; 15'd1753: duty=112; 15'd1754: duty=117; 15'd1755: duty=119; 15'd1756: duty=104; 15'd1757: duty=105; 15'd1758: duty=113; 15'd1759: duty=110;
15'd1760: duty=121; 15'd1761: duty=108; 15'd1762: duty=94; 15'd1763: duty=96; 15'd1764: duty=109; 15'd1765: duty=113; 15'd1766: duty=123; 15'd1767: duty=122;
15'd1768: duty=116; 15'd1769: duty=112; 15'd1770: duty=118; 15'd1771: duty=118; 15'd1772: duty=128; 15'd1773: duty=131; 15'd1774: duty=113; 15'd1775: duty=112;
15'd1776: duty=124; 15'd1777: duty=127; 15'd1778: duty=124; 15'd1779: duty=124; 15'd1780: duty=122; 15'd1781: duty=115; 15'd1782: duty=143; 15'd1783: duty=167;
15'd1784: duty=143; 15'd1785: duty=147; 15'd1786: duty=150; 15'd1787: duty=145; 15'd1788: duty=158; 15'd1789: duty=158; 15'd1790: duty=169; 15'd1791: duty=173;
15'd1792: duty=150; 15'd1793: duty=167; 15'd1794: duty=172; 15'd1795: duty=174; 15'd1796: duty=144; 15'd1797: duty=131; 15'd1798: duty=135; 15'd1799: duty=136;
15'd1800: duty=150; 15'd1801: duty=146; 15'd1802: duty=148; 15'd1803: duty=144; 15'd1804: duty=132; 15'd1805: duty=122; 15'd1806: duty=121; 15'd1807: duty=128;
15'd1808: duty=149; 15'd1809: duty=133; 15'd1810: duty=122; 15'd1811: duty=119; 15'd1812: duty=114; 15'd1813: duty=122; 15'd1814: duty=102; 15'd1815: duty=94;
15'd1816: duty=103; 15'd1817: duty=124; 15'd1818: duty=123; 15'd1819: duty=115; 15'd1820: duty=121; 15'd1821: duty=104; 15'd1822: duty=103; 15'd1823: duty=117;
15'd1824: duty=116; 15'd1825: duty=127; 15'd1826: duty=133; 15'd1827: duty=115; 15'd1828: duty=119; 15'd1829: duty=111; 15'd1830: duty=112; 15'd1831: duty=113;
15'd1832: duty=121; 15'd1833: duty=126; 15'd1834: duty=136; 15'd1835: duty=144; 15'd1836: duty=128; 15'd1837: duty=130; 15'd1838: duty=152; 15'd1839: duty=139;
15'd1840: duty=125; 15'd1841: duty=140; 15'd1842: duty=141; 15'd1843: duty=135; 15'd1844: duty=139; 15'd1845: duty=157; 15'd1846: duty=160; 15'd1847: duty=143;
15'd1848: duty=126; 15'd1849: duty=135; 15'd1850: duty=137; 15'd1851: duty=143; 15'd1852: duty=145; 15'd1853: duty=129; 15'd1854: duty=120; 15'd1855: duty=146;
15'd1856: duty=160; 15'd1857: duty=146; 15'd1858: duty=126; 15'd1859: duty=115; 15'd1860: duty=112; 15'd1861: duty=118; 15'd1862: duty=128; 15'd1863: duty=131;
15'd1864: duty=137; 15'd1865: duty=134; 15'd1866: duty=118; 15'd1867: duty=127; 15'd1868: duty=127; 15'd1869: duty=128; 15'd1870: duty=136; 15'd1871: duty=136;
15'd1872: duty=127; 15'd1873: duty=128; 15'd1874: duty=131; 15'd1875: duty=139; 15'd1876: duty=143; 15'd1877: duty=136; 15'd1878: duty=154; 15'd1879: duty=130;
15'd1880: duty=118; 15'd1881: duty=121; 15'd1882: duty=121; 15'd1883: duty=118; 15'd1884: duty=100; 15'd1885: duty=94; 15'd1886: duty=96; 15'd1887: duty=110;
15'd1888: duty=142; 15'd1889: duty=153; 15'd1890: duty=146; 15'd1891: duty=137; 15'd1892: duty=144; 15'd1893: duty=161; 15'd1894: duty=158; 15'd1895: duty=163;
15'd1896: duty=155; 15'd1897: duty=150; 15'd1898: duty=154; 15'd1899: duty=151; 15'd1900: duty=162; 15'd1901: duty=147; 15'd1902: duty=136; 15'd1903: duty=123;
15'd1904: duty=117; 15'd1905: duty=127; 15'd1906: duty=137; 15'd1907: duty=131; 15'd1908: duty=140; 15'd1909: duty=150; 15'd1910: duty=138; 15'd1911: duty=133;
15'd1912: duty=120; 15'd1913: duty=120; 15'd1914: duty=106; 15'd1915: duty=105; 15'd1916: duty=111; 15'd1917: duty=123; 15'd1918: duty=133; 15'd1919: duty=141;
15'd1920: duty=135; 15'd1921: duty=117; 15'd1922: duty=114; 15'd1923: duty=111; 15'd1924: duty=114; 15'd1925: duty=109; 15'd1926: duty=103; 15'd1927: duty=94;
15'd1928: duty=87; 15'd1929: duty=99; 15'd1930: duty=103; 15'd1931: duty=117; 15'd1932: duty=129; 15'd1933: duty=138; 15'd1934: duty=140; 15'd1935: duty=124;
15'd1936: duty=126; 15'd1937: duty=132; 15'd1938: duty=128; 15'd1939: duty=116; 15'd1940: duty=122; 15'd1941: duty=123; 15'd1942: duty=123; 15'd1943: duty=133;
15'd1944: duty=140; 15'd1945: duty=138; 15'd1946: duty=141; 15'd1947: duty=150; 15'd1948: duty=149; 15'd1949: duty=145; 15'd1950: duty=145; 15'd1951: duty=138;
15'd1952: duty=149; 15'd1953: duty=161; 15'd1954: duty=159; 15'd1955: duty=156; 15'd1956: duty=142; 15'd1957: duty=146; 15'd1958: duty=156; 15'd1959: duty=140;
15'd1960: duty=145; 15'd1961: duty=150; 15'd1962: duty=139; 15'd1963: duty=133; 15'd1964: duty=131; 15'd1965: duty=146; 15'd1966: duty=145; 15'd1967: duty=152;
15'd1968: duty=147; 15'd1969: duty=135; 15'd1970: duty=137; 15'd1971: duty=122; 15'd1972: duty=116; 15'd1973: duty=113; 15'd1974: duty=123; 15'd1975: duty=117;
15'd1976: duty=102; 15'd1977: duty=102; 15'd1978: duty=113; 15'd1979: duty=128; 15'd1980: duty=127; 15'd1981: duty=114; 15'd1982: duty=110; 15'd1983: duty=118;
15'd1984: duty=128; 15'd1985: duty=140; 15'd1986: duty=146; 15'd1987: duty=151; 15'd1988: duty=147; 15'd1989: duty=148; 15'd1990: duty=127; 15'd1991: duty=108;
15'd1992: duty=105; 15'd1993: duty=101; 15'd1994: duty=91; 15'd1995: duty=99; 15'd1996: duty=122; 15'd1997: duty=126; 15'd1998: duty=125; 15'd1999: duty=131;
15'd2000: duty=132; 15'd2001: duty=144; 15'd2002: duty=143; 15'd2003: duty=148; 15'd2004: duty=152; 15'd2005: duty=142; 15'd2006: duty=140; 15'd2007: duty=136;
15'd2008: duty=129; 15'd2009: duty=136; 15'd2010: duty=149; 15'd2011: duty=150; 15'd2012: duty=152; 15'd2013: duty=139; 15'd2014: duty=157; 15'd2015: duty=154;
15'd2016: duty=131; 15'd2017: duty=123; 15'd2018: duty=121; 15'd2019: duty=127; 15'd2020: duty=134; 15'd2021: duty=125; 15'd2022: duty=119; 15'd2023: duty=123;
15'd2024: duty=126; 15'd2025: duty=122; 15'd2026: duty=128; 15'd2027: duty=132; 15'd2028: duty=136; 15'd2029: duty=137; 15'd2030: duty=119; 15'd2031: duty=117;
15'd2032: duty=121; 15'd2033: duty=124; 15'd2034: duty=113; 15'd2035: duty=102; 15'd2036: duty=101; 15'd2037: duty=113; 15'd2038: duty=110; 15'd2039: duty=113;
15'd2040: duty=127; 15'd2041: duty=131; 15'd2042: duty=142; 15'd2043: duty=139; 15'd2044: duty=136; 15'd2045: duty=130; 15'd2046: duty=129; 15'd2047: duty=123;
15'd2048: duty=122; 15'd2049: duty=136; 15'd2050: duty=132; 15'd2051: duty=133; 15'd2052: duty=130; 15'd2053: duty=129; 15'd2054: duty=144; 15'd2055: duty=158;
15'd2056: duty=152; 15'd2057: duty=147; 15'd2058: duty=141; 15'd2059: duty=153; 15'd2060: duty=149; 15'd2061: duty=143; 15'd2062: duty=141; 15'd2063: duty=138;
15'd2064: duty=143; 15'd2065: duty=146; 15'd2066: duty=151; 15'd2067: duty=146; 15'd2068: duty=143; 15'd2069: duty=142; 15'd2070: duty=146; 15'd2071: duty=133;
15'd2072: duty=135; 15'd2073: duty=130; 15'd2074: duty=131; 15'd2075: duty=124; 15'd2076: duty=108; 15'd2077: duty=121; 15'd2078: duty=119; 15'd2079: duty=115;
15'd2080: duty=121; 15'd2081: duty=131; 15'd2082: duty=131; 15'd2083: duty=131; 15'd2084: duty=131; 15'd2085: duty=123; 15'd2086: duty=119; 15'd2087: duty=110;
15'd2088: duty=124; 15'd2089: duty=108; 15'd2090: duty=98; 15'd2091: duty=102; 15'd2092: duty=118; 15'd2093: duty=132; 15'd2094: duty=132; 15'd2095: duty=149;
15'd2096: duty=159; 15'd2097: duty=149; 15'd2098: duty=134; 15'd2099: duty=115; 15'd2100: duty=108; 15'd2101: duty=120; 15'd2102: duty=109; 15'd2103: duty=114;
15'd2104: duty=120; 15'd2105: duty=141; 15'd2106: duty=137; 15'd2107: duty=140; 15'd2108: duty=144; 15'd2109: duty=155; 15'd2110: duty=151; 15'd2111: duty=135;
15'd2112: duty=148; 15'd2113: duty=130; 15'd2114: duty=117; 15'd2115: duty=122; 15'd2116: duty=120; 15'd2117: duty=129; 15'd2118: duty=153; 15'd2119: duty=138;
15'd2120: duty=129; 15'd2121: duty=146; 15'd2122: duty=149; 15'd2123: duty=137; 15'd2124: duty=127; 15'd2125: duty=121; 15'd2126: duty=135; 15'd2127: duty=120;
15'd2128: duty=126; 15'd2129: duty=133; 15'd2130: duty=124; 15'd2131: duty=122; 15'd2132: duty=135; 15'd2133: duty=128; 15'd2134: duty=117; 15'd2135: duty=127;
15'd2136: duty=130; 15'd2137: duty=134; 15'd2138: duty=121; 15'd2139: duty=131; 15'd2140: duty=123; 15'd2141: duty=113; 15'd2142: duty=97; 15'd2143: duty=107;
15'd2144: duty=106; 15'd2145: duty=125; 15'd2146: duty=142; 15'd2147: duty=136; 15'd2148: duty=140; 15'd2149: duty=134; 15'd2150: duty=140; 15'd2151: duty=139;
15'd2152: duty=142; 15'd2153: duty=140; 15'd2154: duty=139; 15'd2155: duty=128; 15'd2156: duty=118; 15'd2157: duty=123; 15'd2158: duty=125; 15'd2159: duty=124;
15'd2160: duty=127; 15'd2161: duty=134; 15'd2162: duty=144; 15'd2163: duty=164; 15'd2164: duty=139; 15'd2165: duty=131; 15'd2166: duty=157; 15'd2167: duty=153;
15'd2168: duty=146; 15'd2169: duty=150; 15'd2170: duty=146; 15'd2171: duty=145; 15'd2172: duty=133; 15'd2173: duty=110; 15'd2174: duty=124; 15'd2175: duty=139;
15'd2176: duty=133; 15'd2177: duty=140; 15'd2178: duty=137; 15'd2179: duty=140; 15'd2180: duty=145; 15'd2181: duty=117; 15'd2182: duty=121; 15'd2183: duty=130;
15'd2184: duty=136; 15'd2185: duty=133; 15'd2186: duty=127; 15'd2187: duty=128; 15'd2188: duty=127; 15'd2189: duty=108; 15'd2190: duty=115; 15'd2191: duty=116;
15'd2192: duty=109; 15'd2193: duty=111; 15'd2194: duty=103; 15'd2195: duty=99; 15'd2196: duty=105; 15'd2197: duty=119; 15'd2198: duty=132; 15'd2199: duty=119;
15'd2200: duty=117; 15'd2201: duty=138; 15'd2202: duty=143; 15'd2203: duty=151; 15'd2204: duty=147; 15'd2205: duty=149; 15'd2206: duty=137; 15'd2207: duty=135;
15'd2208: duty=126; 15'd2209: duty=125; 15'd2210: duty=136; 15'd2211: duty=129; 15'd2212: duty=117; 15'd2213: duty=126; 15'd2214: duty=134; 15'd2215: duty=145;
15'd2216: duty=142; 15'd2217: duty=139; 15'd2218: duty=137; 15'd2219: duty=122; 15'd2220: duty=136; 15'd2221: duty=150; 15'd2222: duty=144; 15'd2223: duty=135;
15'd2224: duty=137; 15'd2225: duty=144; 15'd2226: duty=142; 15'd2227: duty=147; 15'd2228: duty=137; 15'd2229: duty=138; 15'd2230: duty=140; 15'd2231: duty=136;
15'd2232: duty=142; 15'd2233: duty=132; 15'd2234: duty=126; 15'd2235: duty=110; 15'd2236: duty=125; 15'd2237: duty=125; 15'd2238: duty=122; 15'd2239: duty=102;
15'd2240: duty=98; 15'd2241: duty=114; 15'd2242: duty=116; 15'd2243: duty=112; 15'd2244: duty=127; 15'd2245: duty=135; 15'd2246: duty=127; 15'd2247: duty=124;
15'd2248: duty=122; 15'd2249: duty=106; 15'd2250: duty=91; 15'd2251: duty=110; 15'd2252: duty=109; 15'd2253: duty=106; 15'd2254: duty=102; 15'd2255: duty=109;
15'd2256: duty=126; 15'd2257: duty=136; 15'd2258: duty=138; 15'd2259: duty=145; 15'd2260: duty=150; 15'd2261: duty=157; 15'd2262: duty=159; 15'd2263: duty=145;
15'd2264: duty=132; 15'd2265: duty=139; 15'd2266: duty=137; 15'd2267: duty=127; 15'd2268: duty=137; 15'd2269: duty=139; 15'd2270: duty=147; 15'd2271: duty=145;
15'd2272: duty=152; 15'd2273: duty=159; 15'd2274: duty=151; 15'd2275: duty=148; 15'd2276: duty=146; 15'd2277: duty=147; 15'd2278: duty=145; 15'd2279: duty=133;
15'd2280: duty=122; 15'd2281: duty=137; 15'd2282: duty=143; 15'd2283: duty=136; 15'd2284: duty=116; 15'd2285: duty=128; 15'd2286: duty=139; 15'd2287: duty=118;
15'd2288: duty=111; 15'd2289: duty=107; 15'd2290: duty=115; 15'd2291: duty=118; 15'd2292: duty=129; 15'd2293: duty=121; 15'd2294: duty=108; 15'd2295: duty=110;
15'd2296: duty=112; 15'd2297: duty=100; 15'd2298: duty=105; 15'd2299: duty=139; 15'd2300: duty=144; 15'd2301: duty=133; 15'd2302: duty=129; 15'd2303: duty=123;
15'd2304: duty=108; 15'd2305: duty=113; 15'd2306: duty=129; 15'd2307: duty=117; 15'd2308: duty=117; 15'd2309: duty=109; 15'd2310: duty=114; 15'd2311: duty=155;
15'd2312: duty=157; 15'd2313: duty=145; 15'd2314: duty=146; 15'd2315: duty=144; 15'd2316: duty=140; 15'd2317: duty=130; 15'd2318: duty=138; 15'd2319: duty=139;
15'd2320: duty=120; 15'd2321: duty=115; 15'd2322: duty=135; 15'd2323: duty=160; 15'd2324: duty=159; 15'd2325: duty=156; 15'd2326: duty=157; 15'd2327: duty=148;
15'd2328: duty=157; 15'd2329: duty=159; 15'd2330: duty=148; 15'd2331: duty=142; 15'd2332: duty=130; 15'd2333: duty=143; 15'd2334: duty=130; 15'd2335: duty=126;
15'd2336: duty=148; 15'd2337: duty=121; 15'd2338: duty=116; 15'd2339: duty=122; 15'd2340: duty=115; 15'd2341: duty=124; 15'd2342: duty=138; 15'd2343: duty=132;
15'd2344: duty=128; 15'd2345: duty=130; 15'd2346: duty=121; 15'd2347: duty=118; 15'd2348: duty=113; 15'd2349: duty=118; 15'd2350: duty=115; 15'd2351: duty=106;
15'd2352: duty=103; 15'd2353: duty=122; 15'd2354: duty=128; 15'd2355: duty=110; 15'd2356: duty=115; 15'd2357: duty=115; 15'd2358: duty=128; 15'd2359: duty=119;
15'd2360: duty=115; 15'd2361: duty=129; 15'd2362: duty=119; 15'd2363: duty=132; 15'd2364: duty=148; 15'd2365: duty=148; 15'd2366: duty=147; 15'd2367: duty=139;
15'd2368: duty=133; 15'd2369: duty=142; 15'd2370: duty=141; 15'd2371: duty=131; 15'd2372: duty=133; 15'd2373: duty=128; 15'd2374: duty=118; 15'd2375: duty=105;
15'd2376: duty=133; 15'd2377: duty=144; 15'd2378: duty=130; 15'd2379: duty=136; 15'd2380: duty=139; 15'd2381: duty=154; 15'd2382: duty=142; 15'd2383: duty=147;
15'd2384: duty=140; 15'd2385: duty=135; 15'd2386: duty=141; 15'd2387: duty=154; 15'd2388: duty=153; 15'd2389: duty=137; 15'd2390: duty=145; 15'd2391: duty=151;
15'd2392: duty=159; 15'd2393: duty=141; 15'd2394: duty=153; 15'd2395: duty=133; 15'd2396: duty=116; 15'd2397: duty=110; 15'd2398: duty=116; 15'd2399: duty=136;
15'd2400: duty=119; 15'd2401: duty=126; 15'd2402: duty=119; 15'd2403: duty=113; 15'd2404: duty=118; 15'd2405: duty=104; 15'd2406: duty=102; 15'd2407: duty=107;
15'd2408: duty=116; 15'd2409: duty=121; 15'd2410: duty=113; 15'd2411: duty=116; 15'd2412: duty=103; 15'd2413: duty=98; 15'd2414: duty=113; 15'd2415: duty=130;
15'd2416: duty=128; 15'd2417: duty=133; 15'd2418: duty=122; 15'd2419: duty=127; 15'd2420: duty=127; 15'd2421: duty=127; 15'd2422: duty=129; 15'd2423: duty=123;
15'd2424: duty=125; 15'd2425: duty=133; 15'd2426: duty=134; 15'd2427: duty=118; 15'd2428: duty=128; 15'd2429: duty=138; 15'd2430: duty=154; 15'd2431: duty=156;
15'd2432: duty=162; 15'd2433: duty=165; 15'd2434: duty=154; 15'd2435: duty=148; 15'd2436: duty=158; 15'd2437: duty=157; 15'd2438: duty=160; 15'd2439: duty=152;
15'd2440: duty=147; 15'd2441: duty=149; 15'd2442: duty=155; 15'd2443: duty=160; 15'd2444: duty=161; 15'd2445: duty=164; 15'd2446: duty=135; 15'd2447: duty=117;
15'd2448: duty=122; 15'd2449: duty=124; 15'd2450: duty=128; 15'd2451: duty=126; 15'd2452: duty=143; 15'd2453: duty=133; 15'd2454: duty=129; 15'd2455: duty=138;
15'd2456: duty=127; 15'd2457: duty=112; 15'd2458: duty=96; 15'd2459: duty=99; 15'd2460: duty=108; 15'd2461: duty=106; 15'd2462: duty=117; 15'd2463: duty=118;
15'd2464: duty=110; 15'd2465: duty=102; 15'd2466: duty=85; 15'd2467: duty=97; 15'd2468: duty=91; 15'd2469: duty=101; 15'd2470: duty=98; 15'd2471: duty=101;
15'd2472: duty=100; 15'd2473: duty=117; 15'd2474: duty=134; 15'd2475: duty=139; 15'd2476: duty=129; 15'd2477: duty=128; 15'd2478: duty=124; 15'd2479: duty=128;
15'd2480: duty=131; 15'd2481: duty=123; 15'd2482: duty=129; 15'd2483: duty=136; 15'd2484: duty=141; 15'd2485: duty=145; 15'd2486: duty=159; 15'd2487: duty=161;
15'd2488: duty=170; 15'd2489: duty=153; 15'd2490: duty=160; 15'd2491: duty=144; 15'd2492: duty=148; 15'd2493: duty=151; 15'd2494: duty=147; 15'd2495: duty=150;
15'd2496: duty=162; 15'd2497: duty=175; 15'd2498: duty=165; 15'd2499: duty=139; 15'd2500: duty=151; 15'd2501: duty=154; 15'd2502: duty=128; 15'd2503: duty=128;
15'd2504: duty=126; 15'd2505: duty=133; 15'd2506: duty=134; 15'd2507: duty=134; 15'd2508: duty=118; 15'd2509: duty=112; 15'd2510: duty=108; 15'd2511: duty=107;
15'd2512: duty=125; 15'd2513: duty=128; 15'd2514: duty=121; 15'd2515: duty=110; 15'd2516: duty=96; 15'd2517: duty=101; 15'd2518: duty=110; 15'd2519: duty=113;
15'd2520: duty=120; 15'd2521: duty=126; 15'd2522: duty=122; 15'd2523: duty=122; 15'd2524: duty=111; 15'd2525: duty=123; 15'd2526: duty=116; 15'd2527: duty=115;
15'd2528: duty=128; 15'd2529: duty=148; 15'd2530: duty=140; 15'd2531: duty=124; 15'd2532: duty=132; 15'd2533: duty=123; 15'd2534: duty=133; 15'd2535: duty=121;
15'd2536: duty=127; 15'd2537: duty=126; 15'd2538: duty=131; 15'd2539: duty=150; 15'd2540: duty=154; 15'd2541: duty=144; 15'd2542: duty=131; 15'd2543: duty=140;
15'd2544: duty=142; 15'd2545: duty=145; 15'd2546: duty=151; 15'd2547: duty=148; 15'd2548: duty=160; 15'd2549: duty=160; 15'd2550: duty=144; 15'd2551: duty=151;
15'd2552: duty=144; 15'd2553: duty=133; 15'd2554: duty=133; 15'd2555: duty=135; 15'd2556: duty=144; 15'd2557: duty=145; 15'd2558: duty=152; 15'd2559: duty=160;
15'd2560: duty=149; 15'd2561: duty=148; 15'd2562: duty=147; 15'd2563: duty=135; 15'd2564: duty=119; 15'd2565: duty=108; 15'd2566: duty=113; 15'd2567: duty=101;
15'd2568: duty=96; 15'd2569: duty=102; 15'd2570: duty=106; 15'd2571: duty=108; 15'd2572: duty=101; 15'd2573: duty=105; 15'd2574: duty=103; 15'd2575: duty=102;
15'd2576: duty=106; 15'd2577: duty=115; 15'd2578: duty=127; 15'd2579: duty=120; 15'd2580: duty=121; 15'd2581: duty=135; 15'd2582: duty=133; 15'd2583: duty=142;
15'd2584: duty=134; 15'd2585: duty=128; 15'd2586: duty=116; 15'd2587: duty=106; 15'd2588: duty=128; 15'd2589: duty=127; 15'd2590: duty=124; 15'd2591: duty=114;
15'd2592: duty=105; 15'd2593: duty=124; 15'd2594: duty=135; 15'd2595: duty=128; 15'd2596: duty=144; 15'd2597: duty=158; 15'd2598: duty=153; 15'd2599: duty=157;
15'd2600: duty=174; 15'd2601: duty=172; 15'd2602: duty=157; 15'd2603: duty=139; 15'd2604: duty=136; 15'd2605: duty=138; 15'd2606: duty=149; 15'd2607: duty=149;
15'd2608: duty=159; 15'd2609: duty=155; 15'd2610: duty=132; 15'd2611: duty=141; 15'd2612: duty=138; 15'd2613: duty=149; 15'd2614: duty=146; 15'd2615: duty=136;
15'd2616: duty=128; 15'd2617: duty=126; 15'd2618: duty=137; 15'd2619: duty=115; 15'd2620: duty=113; 15'd2621: duty=102; 15'd2622: duty=102; 15'd2623: duty=121;
15'd2624: duty=100; 15'd2625: duty=98; 15'd2626: duty=100; 15'd2627: duty=125; 15'd2628: duty=139; 15'd2629: duty=134; 15'd2630: duty=134; 15'd2631: duty=127;
15'd2632: duty=120; 15'd2633: duty=113; 15'd2634: duty=105; 15'd2635: duty=112; 15'd2636: duty=113; 15'd2637: duty=113; 15'd2638: duty=116; 15'd2639: duty=113;
15'd2640: duty=123; 15'd2641: duty=124; 15'd2642: duty=118; 15'd2643: duty=125; 15'd2644: duty=128; 15'd2645: duty=125; 15'd2646: duty=124; 15'd2647: duty=128;
15'd2648: duty=141; 15'd2649: duty=144; 15'd2650: duty=142; 15'd2651: duty=145; 15'd2652: duty=159; 15'd2653: duty=162; 15'd2654: duty=153; 15'd2655: duty=143;
15'd2656: duty=146; 15'd2657: duty=134; 15'd2658: duty=148; 15'd2659: duty=156; 15'd2660: duty=151; 15'd2661: duty=150; 15'd2662: duty=142; 15'd2663: duty=140;
15'd2664: duty=142; 15'd2665: duty=151; 15'd2666: duty=149; 15'd2667: duty=157; 15'd2668: duty=147; 15'd2669: duty=139; 15'd2670: duty=151; 15'd2671: duty=143;
15'd2672: duty=131; 15'd2673: duty=115; 15'd2674: duty=110; 15'd2675: duty=118; 15'd2676: duty=122; 15'd2677: duty=126; 15'd2678: duty=125; 15'd2679: duty=115;
15'd2680: duty=111; 15'd2681: duty=114; 15'd2682: duty=112; 15'd2683: duty=114; 15'd2684: duty=112; 15'd2685: duty=120; 15'd2686: duty=108; 15'd2687: duty=98;
15'd2688: duty=116; 15'd2689: duty=126; 15'd2690: duty=130; 15'd2691: duty=145; 15'd2692: duty=130; 15'd2693: duty=113; 15'd2694: duty=117; 15'd2695: duty=115;
15'd2696: duty=119; 15'd2697: duty=116; 15'd2698: duty=117; 15'd2699: duty=126; 15'd2700: duty=135; 15'd2701: duty=131; 15'd2702: duty=143; 15'd2703: duty=148;
15'd2704: duty=128; 15'd2705: duty=130; 15'd2706: duty=132; 15'd2707: duty=146; 15'd2708: duty=148; 15'd2709: duty=151; 15'd2710: duty=154; 15'd2711: duty=158;
15'd2712: duty=162; 15'd2713: duty=141; 15'd2714: duty=144; 15'd2715: duty=139; 15'd2716: duty=130; 15'd2717: duty=127; 15'd2718: duty=129; 15'd2719: duty=134;
15'd2720: duty=139; 15'd2721: duty=141; 15'd2722: duty=127; 15'd2723: duty=138; 15'd2724: duty=140; 15'd2725: duty=128; 15'd2726: duty=126; 15'd2727: duty=113;
15'd2728: duty=114; 15'd2729: duty=118; 15'd2730: duty=110; 15'd2731: duty=90; 15'd2732: duty=100; 15'd2733: duty=106; 15'd2734: duty=116; 15'd2735: duty=129;
15'd2736: duty=122; 15'd2737: duty=141; 15'd2738: duty=146; 15'd2739: duty=148; 15'd2740: duty=148; 15'd2741: duty=142; 15'd2742: duty=154; 15'd2743: duty=134;
15'd2744: duty=121; 15'd2745: duty=122; 15'd2746: duty=132; 15'd2747: duty=130; 15'd2748: duty=119; 15'd2749: duty=116; 15'd2750: duty=113; 15'd2751: duty=137;
15'd2752: duty=139; 15'd2753: duty=142; 15'd2754: duty=154; 15'd2755: duty=159; 15'd2756: duty=128; 15'd2757: duty=121; 15'd2758: duty=134; 15'd2759: duty=139;
15'd2760: duty=132; 15'd2761: duty=136; 15'd2762: duty=124; 15'd2763: duty=127; 15'd2764: duty=145; 15'd2765: duty=150; 15'd2766: duty=161; 15'd2767: duty=147;
15'd2768: duty=152; 15'd2769: duty=138; 15'd2770: duty=132; 15'd2771: duty=130; 15'd2772: duty=131; 15'd2773: duty=144; 15'd2774: duty=133; 15'd2775: duty=139;
15'd2776: duty=141; 15'd2777: duty=127; 15'd2778: duty=111; 15'd2779: duty=104; 15'd2780: duty=116; 15'd2781: duty=112; 15'd2782: duty=114; 15'd2783: duty=112;
15'd2784: duty=105; 15'd2785: duty=120; 15'd2786: duty=125; 15'd2787: duty=117; 15'd2788: duty=96; 15'd2789: duty=92; 15'd2790: duty=112; 15'd2791: duty=113;
15'd2792: duty=113; 15'd2793: duty=115; 15'd2794: duty=134; 15'd2795: duty=144; 15'd2796: duty=131; 15'd2797: duty=134; 15'd2798: duty=131; 15'd2799: duty=128;
15'd2800: duty=129; 15'd2801: duty=137; 15'd2802: duty=152; 15'd2803: duty=165; 15'd2804: duty=168; 15'd2805: duty=131; 15'd2806: duty=119; 15'd2807: duty=130;
15'd2808: duty=131; 15'd2809: duty=130; 15'd2810: duty=104; 15'd2811: duty=107; 15'd2812: duty=122; 15'd2813: duty=125; 15'd2814: duty=135; 15'd2815: duty=153;
15'd2816: duty=157; 15'd2817: duty=150; 15'd2818: duty=152; 15'd2819: duty=177; 15'd2820: duty=168; 15'd2821: duty=151; 15'd2822: duty=140; 15'd2823: duty=120;
15'd2824: duty=141; 15'd2825: duty=150; 15'd2826: duty=143; 15'd2827: duty=128; 15'd2828: duty=124; 15'd2829: duty=129; 15'd2830: duty=134; 15'd2831: duty=138;
15'd2832: duty=128; 15'd2833: duty=113; 15'd2834: duty=104; 15'd2835: duty=106; 15'd2836: duty=119; 15'd2837: duty=113; 15'd2838: duty=113; 15'd2839: duty=128;
15'd2840: duty=121; 15'd2841: duty=134; 15'd2842: duty=143; 15'd2843: duty=131; 15'd2844: duty=128; 15'd2845: duty=125; 15'd2846: duty=107; 15'd2847: duty=117;
15'd2848: duty=133; 15'd2849: duty=141; 15'd2850: duty=137; 15'd2851: duty=123; 15'd2852: duty=143; 15'd2853: duty=137; 15'd2854: duty=130; 15'd2855: duty=134;
15'd2856: duty=129; 15'd2857: duty=118; 15'd2858: duty=125; 15'd2859: duty=130; 15'd2860: duty=126; 15'd2861: duty=123; 15'd2862: duty=122; 15'd2863: duty=116;
15'd2864: duty=114; 15'd2865: duty=128; 15'd2866: duty=148; 15'd2867: duty=155; 15'd2868: duty=154; 15'd2869: duty=150; 15'd2870: duty=127; 15'd2871: duty=132;
15'd2872: duty=133; 15'd2873: duty=140; 15'd2874: duty=147; 15'd2875: duty=138; 15'd2876: duty=138; 15'd2877: duty=142; 15'd2878: duty=138; 15'd2879: duty=129;
15'd2880: duty=121; 15'd2881: duty=120; 15'd2882: duty=120; 15'd2883: duty=129; 15'd2884: duty=129; 15'd2885: duty=122; 15'd2886: duty=128; 15'd2887: duty=122;
15'd2888: duty=137; 15'd2889: duty=121; 15'd2890: duty=115; 15'd2891: duty=114; 15'd2892: duty=106; 15'd2893: duty=119; 15'd2894: duty=119; 15'd2895: duty=119;
15'd2896: duty=119; 15'd2897: duty=124; 15'd2898: duty=115; 15'd2899: duty=126; 15'd2900: duty=141; 15'd2901: duty=140; 15'd2902: duty=122; 15'd2903: duty=107;
15'd2904: duty=126; 15'd2905: duty=127; 15'd2906: duty=139; 15'd2907: duty=140; 15'd2908: duty=127; 15'd2909: duty=134; 15'd2910: duty=137; 15'd2911: duty=133;
15'd2912: duty=124; 15'd2913: duty=129; 15'd2914: duty=136; 15'd2915: duty=140; 15'd2916: duty=158; 15'd2917: duty=162; 15'd2918: duty=149; 15'd2919: duty=145;
15'd2920: duty=141; 15'd2921: duty=143; 15'd2922: duty=138; 15'd2923: duty=141; 15'd2924: duty=147; 15'd2925: duty=154; 15'd2926: duty=152; 15'd2927: duty=158;
15'd2928: duty=155; 15'd2929: duty=124; 15'd2930: duty=119; 15'd2931: duty=119; 15'd2932: duty=133; 15'd2933: duty=132; 15'd2934: duty=122; 15'd2935: duty=126;
15'd2936: duty=114; 15'd2937: duty=124; 15'd2938: duty=133; 15'd2939: duty=139; 15'd2940: duty=135; 15'd2941: duty=124; 15'd2942: duty=116; 15'd2943: duty=98;
15'd2944: duty=109; 15'd2945: duty=115; 15'd2946: duty=111; 15'd2947: duty=116; 15'd2948: duty=103; 15'd2949: duty=100; 15'd2950: duty=123; 15'd2951: duty=126;
15'd2952: duty=129; 15'd2953: duty=122; 15'd2954: duty=125; 15'd2955: duty=126; 15'd2956: duty=142; 15'd2957: duty=154; 15'd2958: duty=132; 15'd2959: duty=146;
15'd2960: duty=139; 15'd2961: duty=129; 15'd2962: duty=139; 15'd2963: duty=137; 15'd2964: duty=126; 15'd2965: duty=120; 15'd2966: duty=128; 15'd2967: duty=148;
15'd2968: duty=145; 15'd2969: duty=145; 15'd2970: duty=140; 15'd2971: duty=127; 15'd2972: duty=151; 15'd2973: duty=157; 15'd2974: duty=156; 15'd2975: duty=153;
15'd2976: duty=136; 15'd2977: duty=134; 15'd2978: duty=132; 15'd2979: duty=142; 15'd2980: duty=148; 15'd2981: duty=135; 15'd2982: duty=131; 15'd2983: duty=130;
15'd2984: duty=128; 15'd2985: duty=137; 15'd2986: duty=139; 15'd2987: duty=131; 15'd2988: duty=131; 15'd2989: duty=144; 15'd2990: duty=138; 15'd2991: duty=126;
15'd2992: duty=116; 15'd2993: duty=103; 15'd2994: duty=108; 15'd2995: duty=106; 15'd2996: duty=103; 15'd2997: duty=109; 15'd2998: duty=111; 15'd2999: duty=106;
15'd3000: duty=110; 15'd3001: duty=101; 15'd3002: duty=97; 15'd3003: duty=109; 15'd3004: duty=109; 15'd3005: duty=109; 15'd3006: duty=106; 15'd3007: duty=97;
15'd3008: duty=109; 15'd3009: duty=143; 15'd3010: duty=134; 15'd3011: duty=137; 15'd3012: duty=149; 15'd3013: duty=132; 15'd3014: duty=141; 15'd3015: duty=144;
15'd3016: duty=146; 15'd3017: duty=150; 15'd3018: duty=135; 15'd3019: duty=125; 15'd3020: duty=138; 15'd3021: duty=149; 15'd3022: duty=143; 15'd3023: duty=145;
15'd3024: duty=143; 15'd3025: duty=135; 15'd3026: duty=149; 15'd3027: duty=158; 15'd3028: duty=157; 15'd3029: duty=165; 15'd3030: duty=150; 15'd3031: duty=139;
15'd3032: duty=149; 15'd3033: duty=153; 15'd3034: duty=153; 15'd3035: duty=136; 15'd3036: duty=124; 15'd3037: duty=127; 15'd3038: duty=125; 15'd3039: duty=125;
15'd3040: duty=139; 15'd3041: duty=150; 15'd3042: duty=139; 15'd3043: duty=138; 15'd3044: duty=118; 15'd3045: duty=116; 15'd3046: duty=130; 15'd3047: duty=127;
15'd3048: duty=120; 15'd3049: duty=104; 15'd3050: duty=111; 15'd3051: duty=103; 15'd3052: duty=101; 15'd3053: duty=108; 15'd3054: duty=106; 15'd3055: duty=108;
15'd3056: duty=123; 15'd3057: duty=126; 15'd3058: duty=129; 15'd3059: duty=123; 15'd3060: duty=117; 15'd3061: duty=120; 15'd3062: duty=122; 15'd3063: duty=138;
15'd3064: duty=122; 15'd3065: duty=122; 15'd3066: duty=130; 15'd3067: duty=130; 15'd3068: duty=132; 15'd3069: duty=128; 15'd3070: duty=138; 15'd3071: duty=143;
15'd3072: duty=138; 15'd3073: duty=141; 15'd3074: duty=152; 15'd3075: duty=154; 15'd3076: duty=152; 15'd3077: duty=146; 15'd3078: duty=127; 15'd3079: duty=133;
15'd3080: duty=134; 15'd3081: duty=125; 15'd3082: duty=144; 15'd3083: duty=155; 15'd3084: duty=157; 15'd3085: duty=161; 15'd3086: duty=158; 15'd3087: duty=160;
15'd3088: duty=163; 15'd3089: duty=158; 15'd3090: duty=150; 15'd3091: duty=140; 15'd3092: duty=129; 15'd3093: duty=125; 15'd3094: duty=120; 15'd3095: duty=110;
15'd3096: duty=111; 15'd3097: duty=117; 15'd3098: duty=115; 15'd3099: duty=129; 15'd3100: duty=135; 15'd3101: duty=127; 15'd3102: duty=126; 15'd3103: duty=124;
15'd3104: duty=121; 15'd3105: duty=116; 15'd3106: duty=110; 15'd3107: duty=98; 15'd3108: duty=97; 15'd3109: duty=84; 15'd3110: duty=98; 15'd3111: duty=105;
15'd3112: duty=102; 15'd3113: duty=107; 15'd3114: duty=113; 15'd3115: duty=118; 15'd3116: duty=131; 15'd3117: duty=127; 15'd3118: duty=119; 15'd3119: duty=127;
15'd3120: duty=126; 15'd3121: duty=139; 15'd3122: duty=136; 15'd3123: duty=137; 15'd3124: duty=142; 15'd3125: duty=147; 15'd3126: duty=138; 15'd3127: duty=135;
15'd3128: duty=150; 15'd3129: duty=158; 15'd3130: duty=147; 15'd3131: duty=146; 15'd3132: duty=147; 15'd3133: duty=151; 15'd3134: duty=150; 15'd3135: duty=138;
15'd3136: duty=132; 15'd3137: duty=141; 15'd3138: duty=159; 15'd3139: duty=163; 15'd3140: duty=152; 15'd3141: duty=142; 15'd3142: duty=143; 15'd3143: duty=140;
15'd3144: duty=140; 15'd3145: duty=134; 15'd3146: duty=132; 15'd3147: duty=108; 15'd3148: duty=103; 15'd3149: duty=113; 15'd3150: duty=130; 15'd3151: duty=138;
15'd3152: duty=120; 15'd3153: duty=116; 15'd3154: duty=126; 15'd3155: duty=133; 15'd3156: duty=120; 15'd3157: duty=118; 15'd3158: duty=108; 15'd3159: duty=102;
15'd3160: duty=106; 15'd3161: duty=106; 15'd3162: duty=112; 15'd3163: duty=111; 15'd3164: duty=112; 15'd3165: duty=113; 15'd3166: duty=115; 15'd3167: duty=119;
15'd3168: duty=133; 15'd3169: duty=134; 15'd3170: duty=133; 15'd3171: duty=139; 15'd3172: duty=136; 15'd3173: duty=148; 15'd3174: duty=145; 15'd3175: duty=137;
15'd3176: duty=135; 15'd3177: duty=127; 15'd3178: duty=127; 15'd3179: duty=127; 15'd3180: duty=134; 15'd3181: duty=141; 15'd3182: duty=145; 15'd3183: duty=159;
15'd3184: duty=163; 15'd3185: duty=159; 15'd3186: duty=136; 15'd3187: duty=135; 15'd3188: duty=132; 15'd3189: duty=148; 15'd3190: duty=143; 15'd3191: duty=139;
15'd3192: duty=143; 15'd3193: duty=135; 15'd3194: duty=146; 15'd3195: duty=148; 15'd3196: duty=163; 15'd3197: duty=152; 15'd3198: duty=125; 15'd3199: duty=109;
15'd3200: duty=125; 15'd3201: duty=125; 15'd3202: duty=125; 15'd3203: duty=121; 15'd3204: duty=120; 15'd3205: duty=110; 15'd3206: duty=120; 15'd3207: duty=131;
15'd3208: duty=120; 15'd3209: duty=117; 15'd3210: duty=110; 15'd3211: duty=107; 15'd3212: duty=113; 15'd3213: duty=113; 15'd3214: duty=101; 15'd3215: duty=100;
15'd3216: duty=94; 15'd3217: duty=89; 15'd3218: duty=94; 15'd3219: duty=95; 15'd3220: duty=101; 15'd3221: duty=99; 15'd3222: duty=102; 15'd3223: duty=129;
15'd3224: duty=129; 15'd3225: duty=134; 15'd3226: duty=134; 15'd3227: duty=149; 15'd3228: duty=157; 15'd3229: duty=153; 15'd3230: duty=147; 15'd3231: duty=143;
15'd3232: duty=154; 15'd3233: duty=165; 15'd3234: duty=162; 15'd3235: duty=163; 15'd3236: duty=174; 15'd3237: duty=164; 15'd3238: duty=151; 15'd3239: duty=142;
15'd3240: duty=145; 15'd3241: duty=160; 15'd3242: duty=150; 15'd3243: duty=154; 15'd3244: duty=160; 15'd3245: duty=159; 15'd3246: duty=167; 15'd3247: duty=160;
15'd3248: duty=153; 15'd3249: duty=150; 15'd3250: duty=148; 15'd3251: duty=139; 15'd3252: duty=143; 15'd3253: duty=139; 15'd3254: duty=139; 15'd3255: duty=124;
15'd3256: duty=106; 15'd3257: duty=112; 15'd3258: duty=119; 15'd3259: duty=124; 15'd3260: duty=110; 15'd3261: duty=109; 15'd3262: duty=115; 15'd3263: duty=113;
15'd3264: duty=110; 15'd3265: duty=103; 15'd3266: duty=102; 15'd3267: duty=107; 15'd3268: duty=95; 15'd3269: duty=83; 15'd3270: duty=99; 15'd3271: duty=106;
15'd3272: duty=111; 15'd3273: duty=101; 15'd3274: duty=104; 15'd3275: duty=113; 15'd3276: duty=119; 15'd3277: duty=121; 15'd3278: duty=113; 15'd3279: duty=116;
15'd3280: duty=122; 15'd3281: duty=119; 15'd3282: duty=122; 15'd3283: duty=130; 15'd3284: duty=134; 15'd3285: duty=140; 15'd3286: duty=134; 15'd3287: duty=130;
15'd3288: duty=131; 15'd3289: duty=136; 15'd3290: duty=141; 15'd3291: duty=146; 15'd3292: duty=150; 15'd3293: duty=157; 15'd3294: duty=136; 15'd3295: duty=134;
15'd3296: duty=142; 15'd3297: duty=155; 15'd3298: duty=154; 15'd3299: duty=142; 15'd3300: duty=154; 15'd3301: duty=159; 15'd3302: duty=165; 15'd3303: duty=161;
15'd3304: duty=156; 15'd3305: duty=146; 15'd3306: duty=145; 15'd3307: duty=142; 15'd3308: duty=136; 15'd3309: duty=124; 15'd3310: duty=136; 15'd3311: duty=141;
15'd3312: duty=119; 15'd3313: duty=119; 15'd3314: duty=118; 15'd3315: duty=122; 15'd3316: duty=119; 15'd3317: duty=113; 15'd3318: duty=124; 15'd3319: duty=114;
15'd3320: duty=113; 15'd3321: duty=108; 15'd3322: duty=114; 15'd3323: duty=113; 15'd3324: duty=110; 15'd3325: duty=122; 15'd3326: duty=101; 15'd3327: duty=104;
15'd3328: duty=116; 15'd3329: duty=107; 15'd3330: duty=102; 15'd3331: duty=107; 15'd3332: duty=118; 15'd3333: duty=133; 15'd3334: duty=136; 15'd3335: duty=142;
15'd3336: duty=150; 15'd3337: duty=142; 15'd3338: duty=134; 15'd3339: duty=145; 15'd3340: duty=146; 15'd3341: duty=148; 15'd3342: duty=143; 15'd3343: duty=128;
15'd3344: duty=134; 15'd3345: duty=145; 15'd3346: duty=143; 15'd3347: duty=140; 15'd3348: duty=135; 15'd3349: duty=147; 15'd3350: duty=162; 15'd3351: duty=165;
15'd3352: duty=154; 15'd3353: duty=153; 15'd3354: duty=156; 15'd3355: duty=139; 15'd3356: duty=136; 15'd3357: duty=151; 15'd3358: duty=151; 15'd3359: duty=148;
15'd3360: duty=142; 15'd3361: duty=131; 15'd3362: duty=139; 15'd3363: duty=119; 15'd3364: duty=112; 15'd3365: duty=122; 15'd3366: duty=134; 15'd3367: duty=131;
15'd3368: duty=125; 15'd3369: duty=125; 15'd3370: duty=124; 15'd3371: duty=121; 15'd3372: duty=116; 15'd3373: duty=104; 15'd3374: duty=103; 15'd3375: duty=107;
15'd3376: duty=102; 15'd3377: duty=110; 15'd3378: duty=109; 15'd3379: duty=108; 15'd3380: duty=110; 15'd3381: duty=112; 15'd3382: duty=111; 15'd3383: duty=107;
15'd3384: duty=109; 15'd3385: duty=119; 15'd3386: duty=118; 15'd3387: duty=128; 15'd3388: duty=136; 15'd3389: duty=132; 15'd3390: duty=148; 15'd3391: duty=149;
15'd3392: duty=142; 15'd3393: duty=137; 15'd3394: duty=123; 15'd3395: duty=129; 15'd3396: duty=141; 15'd3397: duty=140; 15'd3398: duty=136; 15'd3399: duty=148;
15'd3400: duty=148; 15'd3401: duty=153; 15'd3402: duty=144; 15'd3403: duty=139; 15'd3404: duty=145; 15'd3405: duty=137; 15'd3406: duty=133; 15'd3407: duty=153;
15'd3408: duty=160; 15'd3409: duty=158; 15'd3410: duty=152; 15'd3411: duty=145; 15'd3412: duty=148; 15'd3413: duty=150; 15'd3414: duty=136; 15'd3415: duty=119;
15'd3416: duty=131; 15'd3417: duty=139; 15'd3418: duty=140; 15'd3419: duty=136; 15'd3420: duty=134; 15'd3421: duty=121; 15'd3422: duty=130; 15'd3423: duty=121;
15'd3424: duty=124; 15'd3425: duty=122; 15'd3426: duty=124; 15'd3427: duty=116; 15'd3428: duty=96; 15'd3429: duty=93; 15'd3430: duty=99; 15'd3431: duty=101;
15'd3432: duty=93; 15'd3433: duty=93; 15'd3434: duty=108; 15'd3435: duty=126; 15'd3436: duty=111; 15'd3437: duty=104; 15'd3438: duty=111; 15'd3439: duty=123;
15'd3440: duty=124; 15'd3441: duty=120; 15'd3442: duty=122; 15'd3443: duty=129; 15'd3444: duty=133; 15'd3445: duty=128; 15'd3446: duty=128; 15'd3447: duty=136;
15'd3448: duty=139; 15'd3449: duty=144; 15'd3450: duty=139; 15'd3451: duty=142; 15'd3452: duty=149; 15'd3453: duty=141; 15'd3454: duty=140; 15'd3455: duty=141;
15'd3456: duty=141; 15'd3457: duty=144; 15'd3458: duty=138; 15'd3459: duty=139; 15'd3460: duty=152; 15'd3461: duty=159; 15'd3462: duty=146; 15'd3463: duty=137;
15'd3464: duty=137; 15'd3465: duty=139; 15'd3466: duty=148; 15'd3467: duty=141; 15'd3468: duty=129; 15'd3469: duty=133; 15'd3470: duty=132; 15'd3471: duty=124;
15'd3472: duty=131; 15'd3473: duty=133; 15'd3474: duty=135; 15'd3475: duty=134; 15'd3476: duty=131; 15'd3477: duty=130; 15'd3478: duty=133; 15'd3479: duty=133;
15'd3480: duty=114; 15'd3481: duty=119; 15'd3482: duty=119; 15'd3483: duty=111; 15'd3484: duty=110; 15'd3485: duty=110; 15'd3486: duty=122; 15'd3487: duty=121;
15'd3488: duty=127; 15'd3489: duty=134; 15'd3490: duty=134; 15'd3491: duty=129; 15'd3492: duty=136; 15'd3493: duty=127; 15'd3494: duty=124; 15'd3495: duty=132;
15'd3496: duty=131; 15'd3497: duty=133; 15'd3498: duty=138; 15'd3499: duty=145; 15'd3500: duty=145; 15'd3501: duty=146; 15'd3502: duty=141; 15'd3503: duty=147;
15'd3504: duty=150; 15'd3505: duty=149; 15'd3506: duty=145; 15'd3507: duty=140; 15'd3508: duty=140; 15'd3509: duty=137; 15'd3510: duty=133; 15'd3511: duty=134;
15'd3512: duty=136; 15'd3513: duty=142; 15'd3514: duty=144; 15'd3515: duty=140; 15'd3516: duty=133; 15'd3517: duty=133; 15'd3518: duty=142; 15'd3519: duty=143;
15'd3520: duty=136; 15'd3521: duty=124; 15'd3522: duty=124; 15'd3523: duty=122; 15'd3524: duty=119; 15'd3525: duty=124; 15'd3526: duty=126; 15'd3527: duty=118;
15'd3528: duty=116; 15'd3529: duty=122; 15'd3530: duty=119; 15'd3531: duty=120; 15'd3532: duty=124; 15'd3533: duty=123; 15'd3534: duty=116; 15'd3535: duty=113;
15'd3536: duty=111; 15'd3537: duty=105; 15'd3538: duty=101; 15'd3539: duty=99; 15'd3540: duty=107; 15'd3541: duty=104; 15'd3542: duty=105; 15'd3543: duty=114;
15'd3544: duty=118; 15'd3545: duty=121; 15'd3546: duty=121; 15'd3547: duty=126; 15'd3548: duty=129; 15'd3549: duty=126; 15'd3550: duty=125; 15'd3551: duty=131;
15'd3552: duty=136; 15'd3553: duty=133; 15'd3554: duty=133; 15'd3555: duty=139; 15'd3556: duty=140; 15'd3557: duty=147; 15'd3558: duty=148; 15'd3559: duty=155;
15'd3560: duty=157; 15'd3561: duty=151; 15'd3562: duty=150; 15'd3563: duty=149; 15'd3564: duty=154; 15'd3565: duty=153; 15'd3566: duty=150; 15'd3567: duty=148;
15'd3568: duty=147; 15'd3569: duty=145; 15'd3570: duty=144; 15'd3571: duty=142; 15'd3572: duty=144; 15'd3573: duty=148; 15'd3574: duty=145; 15'd3575: duty=139;
15'd3576: duty=134; 15'd3577: duty=127; 15'd3578: duty=127; 15'd3579: duty=115; 15'd3580: duty=114; 15'd3581: duty=119; 15'd3582: duty=121; 15'd3583: duty=119;
15'd3584: duty=111; 15'd3585: duty=113; 15'd3586: duty=116; 15'd3587: duty=119; 15'd3588: duty=104; 15'd3589: duty=102; 15'd3590: duty=101; 15'd3591: duty=103;
15'd3592: duty=111; 15'd3593: duty=109; 15'd3594: duty=110; 15'd3595: duty=115; 15'd3596: duty=119; 15'd3597: duty=127; 15'd3598: duty=124; 15'd3599: duty=123;
15'd3600: duty=132; 15'd3601: duty=127; 15'd3602: duty=125; 15'd3603: duty=136; 15'd3604: duty=139; 15'd3605: duty=144; 15'd3606: duty=153; 15'd3607: duty=150;
15'd3608: duty=151; 15'd3609: duty=153; 15'd3610: duty=151; 15'd3611: duty=156; 15'd3612: duty=156; 15'd3613: duty=159; 15'd3614: duty=162; 15'd3615: duty=156;
15'd3616: duty=152; 15'd3617: duty=145; 15'd3618: duty=152; 15'd3619: duty=153; 15'd3620: duty=151; 15'd3621: duty=148; 15'd3622: duty=145; 15'd3623: duty=153;
15'd3624: duty=152; 15'd3625: duty=149; 15'd3626: duty=146; 15'd3627: duty=144; 15'd3628: duty=142; 15'd3629: duty=134; 15'd3630: duty=131; 15'd3631: duty=127;
15'd3632: duty=128; 15'd3633: duty=128; 15'd3634: duty=127; 15'd3635: duty=121; 15'd3636: duty=119; 15'd3637: duty=116; 15'd3638: duty=115; 15'd3639: duty=118;
15'd3640: duty=115; 15'd3641: duty=113; 15'd3642: duty=107; 15'd3643: duty=99; 15'd3644: duty=100; 15'd3645: duty=102; 15'd3646: duty=95; 15'd3647: duty=101;
15'd3648: duty=103; 15'd3649: duty=100; 15'd3650: duty=101; 15'd3651: duty=104; 15'd3652: duty=101; 15'd3653: duty=107; 15'd3654: duty=106; 15'd3655: duty=107;
15'd3656: duty=116; 15'd3657: duty=116; 15'd3658: duty=118; 15'd3659: duty=120; 15'd3660: duty=126; 15'd3661: duty=132; 15'd3662: duty=129; 15'd3663: duty=131;
15'd3664: duty=135; 15'd3665: duty=138; 15'd3666: duty=139; 15'd3667: duty=139; 15'd3668: duty=145; 15'd3669: duty=142; 15'd3670: duty=142; 15'd3671: duty=142;
15'd3672: duty=145; 15'd3673: duty=148; 15'd3674: duty=150; 15'd3675: duty=151; 15'd3676: duty=156; 15'd3677: duty=157; 15'd3678: duty=151; 15'd3679: duty=153;
15'd3680: duty=157; 15'd3681: duty=154; 15'd3682: duty=153; 15'd3683: duty=149; 15'd3684: duty=142; 15'd3685: duty=142; 15'd3686: duty=144; 15'd3687: duty=145;
15'd3688: duty=137; 15'd3689: duty=139; 15'd3690: duty=147; 15'd3691: duty=141; 15'd3692: duty=134; 15'd3693: duty=129; 15'd3694: duty=127; 15'd3695: duty=125;
15'd3696: duty=122; 15'd3697: duty=118; 15'd3698: duty=115; 15'd3699: duty=114; 15'd3700: duty=113; 15'd3701: duty=113; 15'd3702: duty=113; 15'd3703: duty=114;
15'd3704: duty=119; 15'd3705: duty=125; 15'd3706: duty=121; 15'd3707: duty=118; 15'd3708: duty=119; 15'd3709: duty=127; 15'd3710: duty=128; 15'd3711: duty=124;
15'd3712: duty=127; 15'd3713: duty=132; 15'd3714: duty=133; 15'd3715: duty=134; 15'd3716: duty=128; 15'd3717: duty=128; 15'd3718: duty=131; 15'd3719: duty=131;
15'd3720: duty=135; 15'd3721: duty=139; 15'd3722: duty=144; 15'd3723: duty=146; 15'd3724: duty=145; 15'd3725: duty=138; 15'd3726: duty=133; 15'd3727: duty=135;
15'd3728: duty=134; 15'd3729: duty=132; 15'd3730: duty=136; 15'd3731: duty=133; 15'd3732: duty=134; 15'd3733: duty=134; 15'd3734: duty=136; 15'd3735: duty=137;
15'd3736: duty=128; 15'd3737: duty=121; 15'd3738: duty=128; 15'd3739: duty=129; 15'd3740: duty=128; 15'd3741: duty=133; 15'd3742: duty=130; 15'd3743: duty=130;
15'd3744: duty=137; 15'd3745: duty=145; 15'd3746: duty=139; 15'd3747: duty=130; 15'd3748: duty=129; 15'd3749: duty=128; 15'd3750: duty=124; 15'd3751: duty=121;
15'd3752: duty=115; 15'd3753: duty=109; 15'd3754: duty=107; 15'd3755: duty=113; 15'd3756: duty=109; 15'd3757: duty=113; 15'd3758: duty=113; 15'd3759: duty=114;
15'd3760: duty=118; 15'd3761: duty=119; 15'd3762: duty=122; 15'd3763: duty=122; 15'd3764: duty=116; 15'd3765: duty=124; 15'd3766: duty=127; 15'd3767: duty=118;
15'd3768: duty=120; 15'd3769: duty=130; 15'd3770: duty=133; 15'd3771: duty=128; 15'd3772: duty=130; 15'd3773: duty=131; 15'd3774: duty=136; 15'd3775: duty=137;
15'd3776: duty=140; 15'd3777: duty=132; 15'd3778: duty=133; 15'd3779: duty=140; 15'd3780: duty=148; 15'd3781: duty=145; 15'd3782: duty=142; 15'd3783: duty=150;
15'd3784: duty=150; 15'd3785: duty=147; 15'd3786: duty=142; 15'd3787: duty=137; 15'd3788: duty=144; 15'd3789: duty=146; 15'd3790: duty=142; 15'd3791: duty=138;
15'd3792: duty=138; 15'd3793: duty=141; 15'd3794: duty=135; 15'd3795: duty=134; 15'd3796: duty=139; 15'd3797: duty=139; 15'd3798: duty=139; 15'd3799: duty=145;
15'd3800: duty=134; 15'd3801: duty=138; 15'd3802: duty=141; 15'd3803: duty=134; 15'd3804: duty=130; 15'd3805: duty=125; 15'd3806: duty=121; 15'd3807: duty=122;
15'd3808: duty=121; 15'd3809: duty=125; 15'd3810: duty=126; 15'd3811: duty=113; 15'd3812: duty=113; 15'd3813: duty=127; 15'd3814: duty=133; 15'd3815: duty=130;
15'd3816: duty=128; 15'd3817: duty=130; 15'd3818: duty=134; 15'd3819: duty=136; 15'd3820: duty=128; 15'd3821: duty=130; 15'd3822: duty=139; 15'd3823: duty=142;
15'd3824: duty=140; 15'd3825: duty=134; 15'd3826: duty=136; 15'd3827: duty=141; 15'd3828: duty=142; 15'd3829: duty=130; 15'd3830: duty=125; 15'd3831: duty=127;
15'd3832: duty=129; 15'd3833: duty=130; 15'd3834: duty=127; 15'd3835: duty=124; 15'd3836: duty=128; 15'd3837: duty=126; 15'd3838: duty=124; 15'd3839: duty=121;
15'd3840: duty=121; 15'd3841: duty=124; 15'd3842: duty=129; 15'd3843: duty=119; 15'd3844: duty=112; 15'd3845: duty=112; 15'd3846: duty=112; 15'd3847: duty=119;
15'd3848: duty=123; 15'd3849: duty=125; 15'd3850: duty=124; 15'd3851: duty=121; 15'd3852: duty=121; 15'd3853: duty=128; 15'd3854: duty=126; 15'd3855: duty=124;
15'd3856: duty=126; 15'd3857: duty=127; 15'd3858: duty=124; 15'd3859: duty=121; 15'd3860: duty=118; 15'd3861: duty=119; 15'd3862: duty=128; 15'd3863: duty=128;
15'd3864: duty=125; 15'd3865: duty=124; 15'd3866: duty=124; 15'd3867: duty=132; 15'd3868: duty=131; 15'd3869: duty=129; 15'd3870: duty=127; 15'd3871: duty=131;
15'd3872: duty=137; 15'd3873: duty=137; 15'd3874: duty=139; 15'd3875: duty=140; 15'd3876: duty=142; 15'd3877: duty=145; 15'd3878: duty=147; 15'd3879: duty=143;
15'd3880: duty=140; 15'd3881: duty=142; 15'd3882: duty=145; 15'd3883: duty=147; 15'd3884: duty=145; 15'd3885: duty=144; 15'd3886: duty=145; 15'd3887: duty=148;
15'd3888: duty=153; 15'd3889: duty=148; 15'd3890: duty=146; 15'd3891: duty=148; 15'd3892: duty=146; 15'd3893: duty=153; 15'd3894: duty=148; 15'd3895: duty=144;
15'd3896: duty=146; 15'd3897: duty=145; 15'd3898: duty=139; 15'd3899: duty=134; 15'd3900: duty=128; 15'd3901: duty=128; 15'd3902: duty=137; 15'd3903: duty=134;
15'd3904: duty=131; 15'd3905: duty=128; 15'd3906: duty=137; 15'd3907: duty=130; 15'd3908: duty=125; 15'd3909: duty=121; 15'd3910: duty=116; 15'd3911: duty=112;
15'd3912: duty=110; 15'd3913: duty=103; 15'd3914: duty=101; 15'd3915: duty=101; 15'd3916: duty=101; 15'd3917: duty=101; 15'd3918: duty=96; 15'd3919: duty=100;
15'd3920: duty=101; 15'd3921: duty=104; 15'd3922: duty=107; 15'd3923: duty=113; 15'd3924: duty=115; 15'd3925: duty=104; 15'd3926: duty=101; 15'd3927: duty=112;
15'd3928: duty=114; 15'd3929: duty=116; 15'd3930: duty=128; 15'd3931: duty=134; 15'd3932: duty=138; 15'd3933: duty=142; 15'd3934: duty=137; 15'd3935: duty=142;
15'd3936: duty=140; 15'd3937: duty=145; 15'd3938: duty=143; 15'd3939: duty=139; 15'd3940: duty=140; 15'd3941: duty=150; 15'd3942: duty=154; 15'd3943: duty=147;
15'd3944: duty=152; 15'd3945: duty=154; 15'd3946: duty=154; 15'd3947: duty=158; 15'd3948: duty=154; 15'd3949: duty=151; 15'd3950: duty=149; 15'd3951: duty=147;
15'd3952: duty=143; 15'd3953: duty=141; 15'd3954: duty=146; 15'd3955: duty=145; 15'd3956: duty=142; 15'd3957: duty=141; 15'd3958: duty=143; 15'd3959: duty=144;
15'd3960: duty=148; 15'd3961: duty=140; 15'd3962: duty=133; 15'd3963: duty=134; 15'd3964: duty=129; 15'd3965: duty=124; 15'd3966: duty=118; 15'd3967: duty=110;
15'd3968: duty=115; 15'd3969: duty=115; 15'd3970: duty=113; 15'd3971: duty=116; 15'd3972: duty=111; 15'd3973: duty=107; 15'd3974: duty=104; 15'd3975: duty=107;
15'd3976: duty=110; 15'd3977: duty=109; 15'd3978: duty=107; 15'd3979: duty=109; 15'd3980: duty=113; 15'd3981: duty=118; 15'd3982: duty=116; 15'd3983: duty=112;
15'd3984: duty=113; 15'd3985: duty=124; 15'd3986: duty=119; 15'd3987: duty=118; 15'd3988: duty=121; 15'd3989: duty=122; 15'd3990: duty=127; 15'd3991: duty=128;
15'd3992: duty=133; 15'd3993: duty=134; 15'd3994: duty=140; 15'd3995: duty=151; 15'd3996: duty=154; 15'd3997: duty=153; 15'd3998: duty=156; 15'd3999: duty=156;
15'd4000: duty=153; 15'd4001: duty=154; 15'd4002: duty=160; 15'd4003: duty=151; 15'd4004: duty=150; 15'd4005: duty=150; 15'd4006: duty=143; 15'd4007: duty=148;
15'd4008: duty=151; 15'd4009: duty=143; 15'd4010: duty=150; 15'd4011: duty=151; 15'd4012: duty=151; 15'd4013: duty=157; 15'd4014: duty=153; 15'd4015: duty=149;
15'd4016: duty=146; 15'd4017: duty=146; 15'd4018: duty=140; 15'd4019: duty=134; 15'd4020: duty=130; 15'd4021: duty=124; 15'd4022: duty=122; 15'd4023: duty=121;
15'd4024: duty=118; 15'd4025: duty=122; 15'd4026: duty=119; 15'd4027: duty=116; 15'd4028: duty=114; 15'd4029: duty=115; 15'd4030: duty=108; 15'd4031: duty=100;
15'd4032: duty=105; 15'd4033: duty=107; 15'd4034: duty=108; 15'd4035: duty=107; 15'd4036: duty=101; 15'd4037: duty=104; 15'd4038: duty=113; 15'd4039: duty=118;
15'd4040: duty=118; 15'd4041: duty=116; 15'd4042: duty=119; 15'd4043: duty=121; 15'd4044: duty=122; 15'd4045: duty=119; 15'd4046: duty=116; 15'd4047: duty=121;
15'd4048: duty=124; 15'd4049: duty=126; 15'd4050: duty=131; 15'd4051: duty=133; 15'd4052: duty=137; 15'd4053: duty=137; 15'd4054: duty=139; 15'd4055: duty=142;
15'd4056: duty=140; 15'd4057: duty=140; 15'd4058: duty=133; 15'd4059: duty=136; 15'd4060: duty=134; 15'd4061: duty=140; 15'd4062: duty=139; 15'd4063: duty=140;
15'd4064: duty=142; 15'd4065: duty=145; 15'd4066: duty=151; 15'd4067: duty=151; 15'd4068: duty=151; 15'd4069: duty=147; 15'd4070: duty=156; 15'd4071: duty=148;
15'd4072: duty=138; 15'd4073: duty=134; 15'd4074: duty=136; 15'd4075: duty=133; 15'd4076: duty=133; 15'd4077: duty=134; 15'd4078: duty=133; 15'd4079: duty=131;
15'd4080: duty=128; 15'd4081: duty=128; 15'd4082: duty=128; 15'd4083: duty=125; 15'd4084: duty=119; 15'd4085: duty=115; 15'd4086: duty=107; 15'd4087: duty=115;
15'd4088: duty=115; 15'd4089: duty=110; 15'd4090: duty=107; 15'd4091: duty=110; 15'd4092: duty=119; 15'd4093: duty=121; 15'd4094: duty=121; 15'd4095: duty=118;
15'd4096: duty=124; 15'd4097: duty=128; 15'd4098: duty=128; 15'd4099: duty=126; 15'd4100: duty=129; 15'd4101: duty=136; 15'd4102: duty=136; 15'd4103: duty=134;
15'd4104: duty=131; 15'd4105: duty=136; 15'd4106: duty=139; 15'd4107: duty=140; 15'd4108: duty=139; 15'd4109: duty=144; 15'd4110: duty=148; 15'd4111: duty=142;
15'd4112: duty=139; 15'd4113: duty=147; 15'd4114: duty=154; 15'd4115: duty=150; 15'd4116: duty=149; 15'd4117: duty=150; 15'd4118: duty=148; 15'd4119: duty=152;
15'd4120: duty=156; 15'd4121: duty=154; 15'd4122: duty=151; 15'd4123: duty=150; 15'd4124: duty=145; 15'd4125: duty=137; 15'd4126: duty=142; 15'd4127: duty=143;
15'd4128: duty=134; 15'd4129: duty=128; 15'd4130: duty=131; 15'd4131: duty=127; 15'd4132: duty=127; 15'd4133: duty=131; 15'd4134: duty=124; 15'd4135: duty=122;
15'd4136: duty=124; 15'd4137: duty=122; 15'd4138: duty=116; 15'd4139: duty=110; 15'd4140: duty=102; 15'd4141: duty=102; 15'd4142: duty=101; 15'd4143: duty=98;
15'd4144: duty=96; 15'd4145: duty=105; 15'd4146: duty=109; 15'd4147: duty=111; 15'd4148: duty=108; 15'd4149: duty=102; 15'd4150: duty=111; 15'd4151: duty=116;
15'd4152: duty=110; 15'd4153: duty=113; 15'd4154: duty=118; 15'd4155: duty=119; 15'd4156: duty=123; 15'd4157: duty=122; 15'd4158: duty=127; 15'd4159: duty=127;
15'd4160: duty=131; 15'd4161: duty=135; 15'd4162: duty=139; 15'd4163: duty=147; 15'd4164: duty=141; 15'd4165: duty=134; 15'd4166: duty=136; 15'd4167: duty=136;
15'd4168: duty=137; 15'd4169: duty=134; 15'd4170: duty=134; 15'd4171: duty=134; 15'd4172: duty=144; 15'd4173: duty=150; 15'd4174: duty=145; 15'd4175: duty=148;
15'd4176: duty=157; 15'd4177: duty=164; 15'd4178: duty=157; 15'd4179: duty=154; 15'd4180: duty=154; 15'd4181: duty=157; 15'd4182: duty=151; 15'd4183: duty=145;
15'd4184: duty=140; 15'd4185: duty=139; 15'd4186: duty=145; 15'd4187: duty=145; 15'd4188: duty=142; 15'd4189: duty=134; 15'd4190: duty=139; 15'd4191: duty=142;
15'd4192: duty=133; 15'd4193: duty=133; 15'd4194: duty=127; 15'd4195: duty=119; 15'd4196: duty=115; 15'd4197: duty=112; 15'd4198: duty=114; 15'd4199: duty=109;
15'd4200: duty=108; 15'd4201: duty=109; 15'd4202: duty=108; 15'd4203: duty=107; 15'd4204: duty=110; 15'd4205: duty=106; 15'd4206: duty=104; 15'd4207: duty=104;
15'd4208: duty=107; 15'd4209: duty=104; 15'd4210: duty=107; 15'd4211: duty=112; 15'd4212: duty=121; 15'd4213: duty=121; 15'd4214: duty=123; 15'd4215: duty=128;
15'd4216: duty=131; 15'd4217: duty=139; 15'd4218: duty=139; 15'd4219: duty=143; 15'd4220: duty=139; 15'd4221: duty=142; 15'd4222: duty=143; 15'd4223: duty=143;
15'd4224: duty=140; 15'd4225: duty=142; 15'd4226: duty=142; 15'd4227: duty=139; 15'd4228: duty=147; 15'd4229: duty=145; 15'd4230: duty=151; 15'd4231: duty=159;
15'd4232: duty=154; 15'd4233: duty=154; 15'd4234: duty=149; 15'd4235: duty=151; 15'd4236: duty=150; 15'd4237: duty=146; 15'd4238: duty=143; 15'd4239: duty=147;
15'd4240: duty=142; 15'd4241: duty=140; 15'd4242: duty=136; 15'd4243: duty=130; 15'd4244: duty=128; 15'd4245: duty=137; 15'd4246: duty=137; 15'd4247: duty=130;
15'd4248: duty=131; 15'd4249: duty=125; 15'd4250: duty=125; 15'd4251: duty=116; 15'd4252: duty=111; 15'd4253: duty=110; 15'd4254: duty=107; 15'd4255: duty=104;
15'd4256: duty=113; 15'd4257: duty=115; 15'd4258: duty=116; 15'd4259: duty=115; 15'd4260: duty=114; 15'd4261: duty=115; 15'd4262: duty=113; 15'd4263: duty=106;
15'd4264: duty=108; 15'd4265: duty=113; 15'd4266: duty=121; 15'd4267: duty=123; 15'd4268: duty=122; 15'd4269: duty=122; 15'd4270: duty=125; 15'd4271: duty=131;
15'd4272: duty=132; 15'd4273: duty=136; 15'd4274: duty=134; 15'd4275: duty=133; 15'd4276: duty=131; 15'd4277: duty=130; 15'd4278: duty=131; 15'd4279: duty=131;
15'd4280: duty=134; 15'd4281: duty=130; 15'd4282: duty=125; 15'd4283: duty=133; 15'd4284: duty=137; 15'd4285: duty=141; 15'd4286: duty=140; 15'd4287: duty=151;
15'd4288: duty=158; 15'd4289: duty=156; 15'd4290: duty=149; 15'd4291: duty=142; 15'd4292: duty=148; 15'd4293: duty=151; 15'd4294: duty=143; 15'd4295: duty=147;
15'd4296: duty=149; 15'd4297: duty=153; 15'd4298: duty=149; 15'd4299: duty=139; 15'd4300: duty=129; 15'd4301: duty=134; 15'd4302: duty=139; 15'd4303: duty=133;
15'd4304: duty=131; 15'd4305: duty=127; 15'd4306: duty=127; 15'd4307: duty=124; 15'd4308: duty=125; 15'd4309: duty=119; 15'd4310: duty=122; 15'd4311: duty=122;
15'd4312: duty=118; 15'd4313: duty=121; 15'd4314: duty=122; 15'd4315: duty=122; 15'd4316: duty=118; 15'd4317: duty=113; 15'd4318: duty=116; 15'd4319: duty=116;
15'd4320: duty=115; 15'd4321: duty=119; 15'd4322: duty=123; 15'd4323: duty=122; 15'd4324: duty=124; 15'd4325: duty=125; 15'd4326: duty=127; 15'd4327: duty=125;
15'd4328: duty=127; 15'd4329: duty=128; 15'd4330: duty=131; 15'd4331: duty=131; 15'd4332: duty=127; 15'd4333: duty=127; 15'd4334: duty=127; 15'd4335: duty=134;
15'd4336: duty=134; 15'd4337: duty=133; 15'd4338: duty=137; 15'd4339: duty=142; 15'd4340: duty=147; 15'd4341: duty=147; 15'd4342: duty=145; 15'd4343: duty=148;
15'd4344: duty=143; 15'd4345: duty=144; 15'd4346: duty=142; 15'd4347: duty=139; 15'd4348: duty=137; 15'd4349: duty=141; 15'd4350: duty=142; 15'd4351: duty=137;
15'd4352: duty=135; 15'd4353: duty=136; 15'd4354: duty=131; 15'd4355: duty=128; 15'd4356: duty=132; 15'd4357: duty=130; 15'd4358: duty=128; 15'd4359: duty=128;
15'd4360: duty=127; 15'd4361: duty=126; 15'd4362: duty=122; 15'd4363: duty=124; 15'd4364: duty=127; 15'd4365: duty=131; 15'd4366: duty=127; 15'd4367: duty=120;
15'd4368: duty=119; 15'd4369: duty=116; 15'd4370: duty=116; 15'd4371: duty=115; 15'd4372: duty=116; 15'd4373: duty=117; 15'd4374: duty=121; 15'd4375: duty=117;
15'd4376: duty=122; 15'd4377: duty=131; 15'd4378: duty=128; 15'd4379: duty=125; 15'd4380: duty=127; 15'd4381: duty=128; 15'd4382: duty=132; 15'd4383: duty=135;
15'd4384: duty=131; 15'd4385: duty=127; 15'd4386: duty=127; 15'd4387: duty=132; 15'd4388: duty=131; 15'd4389: duty=132; 15'd4390: duty=133; 15'd4391: duty=128;
15'd4392: duty=129; 15'd4393: duty=132; 15'd4394: duty=127; 15'd4395: duty=129; 15'd4396: duty=133; 15'd4397: duty=135; 15'd4398: duty=138; 15'd4399: duty=146;
15'd4400: duty=152; 15'd4401: duty=154; 15'd4402: duty=156; 15'd4403: duty=151; 15'd4404: duty=147; 15'd4405: duty=143; 15'd4406: duty=145; 15'd4407: duty=142;
15'd4408: duty=136; 15'd4409: duty=140; 15'd4410: duty=145; 15'd4411: duty=137; 15'd4412: duty=127; 15'd4413: duty=125; 15'd4414: duty=128; 15'd4415: duty=137;
15'd4416: duty=136; 15'd4417: duty=134; 15'd4418: duty=131; 15'd4419: duty=130; 15'd4420: duty=129; 15'd4421: duty=127; 15'd4422: duty=125; 15'd4423: duty=121;
15'd4424: duty=119; 15'd4425: duty=119; 15'd4426: duty=114; 15'd4427: duty=110; 15'd4428: duty=114; 15'd4429: duty=110; 15'd4430: duty=111; 15'd4431: duty=116;
15'd4432: duty=117; 15'd4433: duty=124; 15'd4434: duty=127; 15'd4435: duty=124; 15'd4436: duty=127; 15'd4437: duty=126; 15'd4438: duty=125; 15'd4439: duty=126;
15'd4440: duty=131; 15'd4441: duty=134; 15'd4442: duty=133; 15'd4443: duty=136; 15'd4444: duty=134; 15'd4445: duty=134; 15'd4446: duty=137; 15'd4447: duty=144;
15'd4448: duty=142; 15'd4449: duty=136; 15'd4450: duty=142; 15'd4451: duty=136; 15'd4452: duty=136; 15'd4453: duty=131; 15'd4454: duty=134; 15'd4455: duty=140;
15'd4456: duty=141; 15'd4457: duty=142; 15'd4458: duty=142; 15'd4459: duty=140; 15'd4460: duty=134; 15'd4461: duty=143; 15'd4462: duty=145; 15'd4463: duty=135;
15'd4464: duty=136; 15'd4465: duty=134; 15'd4466: duty=134; 15'd4467: duty=128; 15'd4468: duty=124; 15'd4469: duty=131; 15'd4470: duty=131; 15'd4471: duty=134;
15'd4472: duty=127; 15'd4473: duty=124; 15'd4474: duty=127; 15'd4475: duty=124; 15'd4476: duty=121; 15'd4477: duty=122; 15'd4478: duty=120; 15'd4479: duty=122;
15'd4480: duty=118; 15'd4481: duty=113; 15'd4482: duty=118; 15'd4483: duty=116; 15'd4484: duty=119; 15'd4485: duty=124; 15'd4486: duty=123; 15'd4487: duty=126;
15'd4488: duty=128; 15'd4489: duty=127; 15'd4490: duty=125; 15'd4491: duty=128; 15'd4492: duty=134; 15'd4493: duty=130; 15'd4494: duty=124; 15'd4495: duty=130;
15'd4496: duty=137; 15'd4497: duty=131; 15'd4498: duty=130; 15'd4499: duty=131; 15'd4500: duty=130; 15'd4501: duty=130; 15'd4502: duty=131; 15'd4503: duty=127;
15'd4504: duty=125; 15'd4505: duty=126; 15'd4506: duty=121; 15'd4507: duty=124; 15'd4508: duty=128; 15'd4509: duty=127; 15'd4510: duty=132; 15'd4511: duty=140;
15'd4512: duty=137; 15'd4513: duty=140; 15'd4514: duty=150; 15'd4515: duty=147; 15'd4516: duty=137; 15'd4517: duty=136; 15'd4518: duty=140; 15'd4519: duty=140;
15'd4520: duty=137; 15'd4521: duty=140; 15'd4522: duty=146; 15'd4523: duty=145; 15'd4524: duty=137; 15'd4525: duty=139; 15'd4526: duty=139; 15'd4527: duty=134;
15'd4528: duty=129; 15'd4529: duty=131; 15'd4530: duty=131; 15'd4531: duty=125; 15'd4532: duty=124; 15'd4533: duty=128; 15'd4534: duty=127; 15'd4535: duty=125;
15'd4536: duty=128; 15'd4537: duty=128; 15'd4538: duty=129; 15'd4539: duty=124; 15'd4540: duty=122; 15'd4541: duty=118; 15'd4542: duty=118; 15'd4543: duty=122;
15'd4544: duty=121; 15'd4545: duty=128; 15'd4546: duty=130; 15'd4547: duty=129; 15'd4548: duty=130; 15'd4549: duty=132; 15'd4550: duty=131; 15'd4551: duty=131;
15'd4552: duty=136; 15'd4553: duty=132; 15'd4554: duty=130; 15'd4555: duty=131; 15'd4556: duty=136; 15'd4557: duty=137; 15'd4558: duty=131; 15'd4559: duty=134;
15'd4560: duty=137; 15'd4561: duty=133; 15'd4562: duty=136; 15'd4563: duty=137; 15'd4564: duty=140; 15'd4565: duty=132; 15'd4566: duty=134; 15'd4567: duty=140;
15'd4568: duty=136; 15'd4569: duty=142; 15'd4570: duty=143; 15'd4571: duty=134; 15'd4572: duty=133; 15'd4573: duty=131; 15'd4574: duty=130; 15'd4575: duty=132;
15'd4576: duty=129; 15'd4577: duty=132; 15'd4578: duty=136; 15'd4579: duty=134; 15'd4580: duty=130; 15'd4581: duty=128; 15'd4582: duty=125; 15'd4583: duty=131;
15'd4584: duty=131; 15'd4585: duty=122; 15'd4586: duty=119; 15'd4587: duty=113; 15'd4588: duty=113; 15'd4589: duty=121; 15'd4590: duty=118; 15'd4591: duty=118;
15'd4592: duty=121; 15'd4593: duty=118; 15'd4594: duty=119; 15'd4595: duty=118; 15'd4596: duty=112; 15'd4597: duty=113; 15'd4598: duty=119; 15'd4599: duty=122;
15'd4600: duty=124; 15'd4601: duty=126; 15'd4602: duty=129; 15'd4603: duty=130; 15'd4604: duty=131; 15'd4605: duty=133; 15'd4606: duty=133; 15'd4607: duty=131;
15'd4608: duty=129; 15'd4609: duty=131; 15'd4610: duty=136; 15'd4611: duty=137; 15'd4612: duty=142; 15'd4613: duty=144; 15'd4614: duty=142; 15'd4615: duty=137;
15'd4616: duty=140; 15'd4617: duty=144; 15'd4618: duty=139; 15'd4619: duty=131; 15'd4620: duty=136; 15'd4621: duty=142; 15'd4622: duty=139; 15'd4623: duty=137;
15'd4624: duty=142; 15'd4625: duty=142; 15'd4626: duty=137; 15'd4627: duty=145; 15'd4628: duty=151; 15'd4629: duty=147; 15'd4630: duty=142; 15'd4631: duty=142;
15'd4632: duty=140; 15'd4633: duty=136; 15'd4634: duty=134; 15'd4635: duty=134; 15'd4636: duty=133; 15'd4637: duty=136; 15'd4638: duty=137; 15'd4639: duty=136;
15'd4640: duty=133; 15'd4641: duty=134; 15'd4642: duty=134; 15'd4643: duty=137; 15'd4644: duty=128; 15'd4645: duty=121; 15'd4646: duty=119; 15'd4647: duty=120;
15'd4648: duty=118; 15'd4649: duty=116; 15'd4650: duty=114; 15'd4651: duty=115; 15'd4652: duty=113; 15'd4653: duty=107; 15'd4654: duty=110; 15'd4655: duty=110;
15'd4656: duty=118; 15'd4657: duty=122; 15'd4658: duty=124; 15'd4659: duty=121; 15'd4660: duty=119; 15'd4661: duty=125; 15'd4662: duty=129; 15'd4663: duty=125;
15'd4664: duty=125; 15'd4665: duty=130; 15'd4666: duty=134; 15'd4667: duty=137; 15'd4668: duty=140; 15'd4669: duty=140; 15'd4670: duty=137; 15'd4671: duty=133;
15'd4672: duty=130; 15'd4673: duty=134; 15'd4674: duty=139; 15'd4675: duty=140; 15'd4676: duty=143; 15'd4677: duty=143; 15'd4678: duty=144; 15'd4679: duty=146;
15'd4680: duty=142; 15'd4681: duty=137; 15'd4682: duty=134; 15'd4683: duty=136; 15'd4684: duty=142; 15'd4685: duty=134; 15'd4686: duty=129; 15'd4687: duty=133;
15'd4688: duty=139; 15'd4689: duty=139; 15'd4690: duty=131; 15'd4691: duty=130; 15'd4692: duty=131; 15'd4693: duty=133; 15'd4694: duty=129; 15'd4695: duty=124;
15'd4696: duty=121; 15'd4697: duty=129; 15'd4698: duty=128; 15'd4699: duty=121; 15'd4700: duty=116; 15'd4701: duty=116; 15'd4702: duty=124; 15'd4703: duty=125;
15'd4704: duty=125; 15'd4705: duty=124; 15'd4706: duty=122; 15'd4707: duty=119; 15'd4708: duty=115; 15'd4709: duty=109; 15'd4710: duty=108; 15'd4711: duty=115;
15'd4712: duty=122; 15'd4713: duty=122; 15'd4714: duty=125; 15'd4715: duty=126; 15'd4716: duty=128; 15'd4717: duty=131; 15'd4718: duty=132; 15'd4719: duty=131;
15'd4720: duty=131; 15'd4721: duty=134; 15'd4722: duty=134; 15'd4723: duty=134; 15'd4724: duty=134; 15'd4725: duty=142; 15'd4726: duty=148; 15'd4727: duty=144;
15'd4728: duty=148; 15'd4729: duty=153; 15'd4730: duty=149; 15'd4731: duty=145; 15'd4732: duty=137; 15'd4733: duty=136; 15'd4734: duty=137; 15'd4735: duty=142;
15'd4736: duty=137; 15'd4737: duty=129; 15'd4738: duty=139; 15'd4739: duty=146; 15'd4740: duty=143; 15'd4741: duty=143; 15'd4742: duty=145; 15'd4743: duty=145;
15'd4744: duty=147; 15'd4745: duty=142; 15'd4746: duty=137; 15'd4747: duty=139; 15'd4748: duty=144; 15'd4749: duty=139; 15'd4750: duty=131; 15'd4751: duty=125;
15'd4752: duty=125; 15'd4753: duty=128; 15'd4754: duty=124; 15'd4755: duty=119; 15'd4756: duty=116; 15'd4757: duty=115; 15'd4758: duty=112; 15'd4759: duty=108;
15'd4760: duty=107; 15'd4761: duty=116; 15'd4762: duty=116; 15'd4763: duty=116; 15'd4764: duty=119; 15'd4765: duty=116; 15'd4766: duty=113; 15'd4767: duty=111;
15'd4768: duty=108; 15'd4769: duty=107; 15'd4770: duty=112; 15'd4771: duty=115; 15'd4772: duty=112; 15'd4773: duty=115; 15'd4774: duty=122; 15'd4775: duty=128;
15'd4776: duty=132; 15'd4777: duty=128; 15'd4778: duty=130; 15'd4779: duty=136; 15'd4780: duty=140; 15'd4781: duty=137; 15'd4782: duty=134; 15'd4783: duty=133;
15'd4784: duty=140; 15'd4785: duty=145; 15'd4786: duty=142; 15'd4787: duty=139; 15'd4788: duty=142; 15'd4789: duty=151; 15'd4790: duty=154; 15'd4791: duty=151;
15'd4792: duty=148; 15'd4793: duty=150; 15'd4794: duty=151; 15'd4795: duty=147; 15'd4796: duty=145; 15'd4797: duty=147; 15'd4798: duty=154; 15'd4799: duty=157;
15'd4800: duty=146; 15'd4801: duty=144; 15'd4802: duty=143; 15'd4803: duty=145; 15'd4804: duty=143; 15'd4805: duty=131; 15'd4806: duty=128; 15'd4807: duty=130;
15'd4808: duty=129; 15'd4809: duty=127; 15'd4810: duty=127; 15'd4811: duty=125; 15'd4812: duty=124; 15'd4813: duty=121; 15'd4814: duty=113; 15'd4815: duty=115;
15'd4816: duty=116; 15'd4817: duty=115; 15'd4818: duty=115; 15'd4819: duty=112; 15'd4820: duty=112; 15'd4821: duty=112; 15'd4822: duty=107; 15'd4823: duty=99;
15'd4824: duty=98; 15'd4825: duty=110; 15'd4826: duty=118; 15'd4827: duty=116; 15'd4828: duty=116; 15'd4829: duty=118; 15'd4830: duty=124; 15'd4831: duty=128;
15'd4832: duty=119; 15'd4833: duty=119; 15'd4834: duty=131; 15'd4835: duty=131; 15'd4836: duty=128; 15'd4837: duty=125; 15'd4838: duty=131; 15'd4839: duty=137;
15'd4840: duty=139; 15'd4841: duty=135; 15'd4842: duty=136; 15'd4843: duty=142; 15'd4844: duty=147; 15'd4845: duty=143; 15'd4846: duty=140; 15'd4847: duty=136;
15'd4848: duty=139; 15'd4849: duty=149; 15'd4850: duty=150; 15'd4851: duty=140; 15'd4852: duty=142; 15'd4853: duty=151; 15'd4854: duty=147; 15'd4855: duty=148;
15'd4856: duty=145; 15'd4857: duty=146; 15'd4858: duty=140; 15'd4859: duty=142; 15'd4860: duty=145; 15'd4861: duty=142; 15'd4862: duty=143; 15'd4863: duty=148;
15'd4864: duty=148; 15'd4865: duty=143; 15'd4866: duty=140; 15'd4867: duty=142; 15'd4868: duty=134; 15'd4869: duty=125; 15'd4870: duty=126; 15'd4871: duty=127;
15'd4872: duty=121; 15'd4873: duty=112; 15'd4874: duty=105; 15'd4875: duty=112; 15'd4876: duty=124; 15'd4877: duty=119; 15'd4878: duty=111; 15'd4879: duty=107;
15'd4880: duty=109; 15'd4881: duty=107; 15'd4882: duty=104; 15'd4883: duty=101; 15'd4884: duty=106; 15'd4885: duty=118; 15'd4886: duty=119; 15'd4887: duty=119;
15'd4888: duty=124; 15'd4889: duty=126; 15'd4890: duty=134; 15'd4891: duty=133; 15'd4892: duty=128; 15'd4893: duty=122; 15'd4894: duty=127; 15'd4895: duty=131;
15'd4896: duty=127; 15'd4897: duty=121; 15'd4898: duty=127; 15'd4899: duty=137; 15'd4900: duty=137; 15'd4901: duty=142; 15'd4902: duty=145; 15'd4903: duty=150;
15'd4904: duty=150; 15'd4905: duty=150; 15'd4906: duty=151; 15'd4907: duty=150; 15'd4908: duty=150; 15'd4909: duty=148; 15'd4910: duty=145; 15'd4911: duty=145;
15'd4912: duty=148; 15'd4913: duty=154; 15'd4914: duty=156; 15'd4915: duty=145; 15'd4916: duty=142; 15'd4917: duty=147; 15'd4918: duty=144; 15'd4919: duty=142;
15'd4920: duty=142; 15'd4921: duty=143; 15'd4922: duty=141; 15'd4923: duty=140; 15'd4924: duty=134; 15'd4925: duty=128; 15'd4926: duty=125; 15'd4927: duty=125;
15'd4928: duty=124; 15'd4929: duty=116; 15'd4930: duty=113; 15'd4931: duty=112; 15'd4932: duty=115; 15'd4933: duty=116; 15'd4934: duty=112; 15'd4935: duty=110;
15'd4936: duty=105; 15'd4937: duty=101; 15'd4938: duty=96; 15'd4939: duty=99; 15'd4940: duty=108; 15'd4941: duty=113; 15'd4942: duty=114; 15'd4943: duty=110;
15'd4944: duty=114; 15'd4945: duty=116; 15'd4946: duty=116; 15'd4947: duty=116; 15'd4948: duty=119; 15'd4949: duty=124; 15'd4950: duty=129; 15'd4951: duty=136;
15'd4952: duty=132; 15'd4953: duty=131; 15'd4954: duty=137; 15'd4955: duty=139; 15'd4956: duty=140; 15'd4957: duty=137; 15'd4958: duty=137; 15'd4959: duty=141;
15'd4960: duty=143; 15'd4961: duty=139; 15'd4962: duty=137; 15'd4963: duty=141; 15'd4964: duty=145; 15'd4965: duty=145; 15'd4966: duty=145; 15'd4967: duty=141;
15'd4968: duty=143; 15'd4969: duty=153; 15'd4970: duty=152; 15'd4971: duty=150; 15'd4972: duty=145; 15'd4973: duty=139; 15'd4974: duty=140; 15'd4975: duty=141;
15'd4976: duty=140; 15'd4977: duty=141; 15'd4978: duty=140; 15'd4979: duty=139; 15'd4980: duty=136; 15'd4981: duty=137; 15'd4982: duty=136; 15'd4983: duty=133;
15'd4984: duty=129; 15'd4985: duty=130; 15'd4986: duty=128; 15'd4987: duty=124; 15'd4988: duty=119; 15'd4989: duty=116; 15'd4990: duty=121; 15'd4991: duty=118;
15'd4992: duty=115; 15'd4993: duty=112; 15'd4994: duty=118; 15'd4995: duty=112; 15'd4996: duty=110; 15'd4997: duty=113; 15'd4998: duty=116; 15'd4999: duty=121;
15'd5000: duty=128; 15'd5001: duty=127; 15'd5002: duty=124; 15'd5003: duty=127; 15'd5004: duty=126; 15'd5005: duty=133; 15'd5006: duty=134; 15'd5007: duty=129;
15'd5008: duty=133; 15'd5009: duty=136; 15'd5010: duty=136; 15'd5011: duty=134; 15'd5012: duty=133; 15'd5013: duty=137; 15'd5014: duty=133; 15'd5015: duty=131;
15'd5016: duty=132; 15'd5017: duty=135; 15'd5018: duty=137; 15'd5019: duty=142; 15'd5020: duty=146; 15'd5021: duty=146; 15'd5022: duty=142; 15'd5023: duty=147;
15'd5024: duty=146; 15'd5025: duty=143; 15'd5026: duty=149; 15'd5027: duty=146; 15'd5028: duty=142; 15'd5029: duty=140; 15'd5030: duty=137; 15'd5031: duty=134;
15'd5032: duty=139; 15'd5033: duty=137; 15'd5034: duty=134; 15'd5035: duty=131; 15'd5036: duty=130; 15'd5037: duty=133; 15'd5038: duty=132; 15'd5039: duty=126;
15'd5040: duty=119; 15'd5041: duty=115; 15'd5042: duty=118; 15'd5043: duty=121; 15'd5044: duty=119; 15'd5045: duty=120; 15'd5046: duty=118; 15'd5047: duty=118;
15'd5048: duty=118; 15'd5049: duty=115; 15'd5050: duty=112; 15'd5051: duty=115; 15'd5052: duty=113; 15'd5053: duty=104; 15'd5054: duty=105; 15'd5055: duty=113;
15'd5056: duty=118; 15'd5057: duty=121; 15'd5058: duty=121; 15'd5059: duty=118; 15'd5060: duty=124; 15'd5061: duty=124; 15'd5062: duty=121; 15'd5063: duty=129;
15'd5064: duty=126; 15'd5065: duty=128; 15'd5066: duty=136; 15'd5067: duty=136; 15'd5068: duty=137; 15'd5069: duty=143; 15'd5070: duty=144; 15'd5071: duty=143;
15'd5072: duty=143; 15'd5073: duty=145; 15'd5074: duty=150; 15'd5075: duty=151; 15'd5076: duty=145; 15'd5077: duty=142; 15'd5078: duty=137; 15'd5079: duty=140;
15'd5080: duty=145; 15'd5081: duty=145; 15'd5082: duty=142; 15'd5083: duty=140; 15'd5084: duty=147; 15'd5085: duty=149; 15'd5086: duty=154; 15'd5087: duty=157;
15'd5088: duty=151; 15'd5089: duty=147; 15'd5090: duty=144; 15'd5091: duty=137; 15'd5092: duty=131; 15'd5093: duty=134; 15'd5094: duty=136; 15'd5095: duty=131;
15'd5096: duty=130; 15'd5097: duty=131; 15'd5098: duty=127; 15'd5099: duty=124; 15'd5100: duty=127; 15'd5101: duty=125; 15'd5102: duty=119; 15'd5103: duty=119;
15'd5104: duty=122; 15'd5105: duty=121; 15'd5106: duty=118; 15'd5107: duty=115; 15'd5108: duty=112; 15'd5109: duty=119; 15'd5110: duty=110; 15'd5111: duty=99;
15'd5112: duty=104; 15'd5113: duty=107; 15'd5114: duty=107; 15'd5115: duty=109; 15'd5116: duty=116; 15'd5117: duty=121; 15'd5118: duty=121; 15'd5119: duty=124;
15'd5120: duty=128; 15'd5121: duty=128; 15'd5122: duty=127; 15'd5123: duty=131; 15'd5124: duty=129; 15'd5125: duty=125; 15'd5126: duty=125; 15'd5127: duty=125;
15'd5128: duty=124; 15'd5129: duty=122; 15'd5130: duty=124; 15'd5131: duty=127; 15'd5132: duty=134; 15'd5133: duty=134; 15'd5134: duty=137; 15'd5135: duty=146;
15'd5136: duty=154; 15'd5137: duty=154; 15'd5138: duty=151; 15'd5139: duty=148; 15'd5140: duty=150; 15'd5141: duty=154; 15'd5142: duty=149; 15'd5143: duty=143;
15'd5144: duty=142; 15'd5145: duty=142; 15'd5146: duty=143; 15'd5147: duty=142; 15'd5148: duty=142; 15'd5149: duty=146; 15'd5150: duty=147; 15'd5151: duty=146;
15'd5152: duty=143; 15'd5153: duty=140; 15'd5154: duty=139; 15'd5155: duty=137; 15'd5156: duty=131; 15'd5157: duty=130; 15'd5158: duty=130; 15'd5159: duty=134;
15'd5160: duty=133; 15'd5161: duty=125; 15'd5162: duty=122; 15'd5163: duty=124; 15'd5164: duty=121; 15'd5165: duty=115; 15'd5166: duty=112; 15'd5167: duty=112;
15'd5168: duty=110; 15'd5169: duty=108; 15'd5170: duty=110; 15'd5171: duty=115; 15'd5172: duty=119; 15'd5173: duty=124; 15'd5174: duty=122; 15'd5175: duty=119;
15'd5176: duty=124; 15'd5177: duty=122; 15'd5178: duty=122; 15'd5179: duty=124; 15'd5180: duty=124; 15'd5181: duty=121; 15'd5182: duty=129; 15'd5183: duty=131;
15'd5184: duty=128; 15'd5185: duty=128; 15'd5186: duty=137; 15'd5187: duty=143; 15'd5188: duty=142; 15'd5189: duty=141; 15'd5190: duty=139; 15'd5191: duty=134;
15'd5192: duty=137; 15'd5193: duty=133; 15'd5194: duty=133; 15'd5195: duty=140; 15'd5196: duty=140; 15'd5197: duty=139; 15'd5198: duty=140; 15'd5199: duty=143;
15'd5200: duty=139; 15'd5201: duty=139; 15'd5202: duty=143; 15'd5203: duty=139; 15'd5204: duty=134; 15'd5205: duty=137; 15'd5206: duty=139; 15'd5207: duty=140;
15'd5208: duty=140; 15'd5209: duty=143; 15'd5210: duty=140; 15'd5211: duty=133; 15'd5212: duty=133; 15'd5213: duty=131; 15'd5214: duty=127; 15'd5215: duty=126;
15'd5216: duty=128; 15'd5217: duty=131; 15'd5218: duty=130; 15'd5219: duty=126; 15'd5220: duty=125; 15'd5221: duty=127; 15'd5222: duty=122; 15'd5223: duty=122;
15'd5224: duty=122; 15'd5225: duty=121; 15'd5226: duty=113; 15'd5227: duty=109; 15'd5228: duty=116; 15'd5229: duty=116; 15'd5230: duty=115; 15'd5231: duty=114;
15'd5232: duty=124; 15'd5233: duty=124; 15'd5234: duty=121; 15'd5235: duty=122; 15'd5236: duty=127; 15'd5237: duty=130; 15'd5238: duty=129; 15'd5239: duty=131;
15'd5240: duty=128; 15'd5241: duty=127; 15'd5242: duty=134; 15'd5243: duty=134; 15'd5244: duty=133; 15'd5245: duty=130; 15'd5246: duty=127; 15'd5247: duty=129;
15'd5248: duty=136; 15'd5249: duty=136; 15'd5250: duty=139; 15'd5251: duty=141; 15'd5252: duty=137; 15'd5253: duty=143; 15'd5254: duty=144; 15'd5255: duty=138;
15'd5256: duty=140; 15'd5257: duty=145; 15'd5258: duty=136; 15'd5259: duty=139; 15'd5260: duty=142; 15'd5261: duty=140; 15'd5262: duty=143; 15'd5263: duty=145;
15'd5264: duty=145; 15'd5265: duty=139; 15'd5266: duty=136; 15'd5267: duty=139; 15'd5268: duty=134; 15'd5269: duty=127; 15'd5270: duty=122; 15'd5271: duty=116;
15'd5272: duty=110; 15'd5273: duty=113; 15'd5274: duty=121; 15'd5275: duty=130; 15'd5276: duty=137; 15'd5277: duty=137; 15'd5278: duty=139; 15'd5279: duty=131;
15'd5280: duty=129; 15'd5281: duty=130; 15'd5282: duty=121; 15'd5283: duty=113; 15'd5284: duty=116; 15'd5285: duty=107; 15'd5286: duty=99; 15'd5287: duty=103;
15'd5288: duty=104; 15'd5289: duty=109; 15'd5290: duty=115; 15'd5291: duty=107; 15'd5292: duty=113; 15'd5293: duty=124; 15'd5294: duty=133; 15'd5295: duty=140;
15'd5296: duty=134; 15'd5297: duty=136; 15'd5298: duty=146; 15'd5299: duty=148; 15'd5300: duty=149; 15'd5301: duty=145; 15'd5302: duty=142; 15'd5303: duty=146;
15'd5304: duty=145; 15'd5305: duty=147; 15'd5306: duty=143; 15'd5307: duty=145; 15'd5308: duty=148; 15'd5309: duty=153; 15'd5310: duty=154; 15'd5311: duty=150;
15'd5312: duty=151; 15'd5313: duty=160; 15'd5314: duty=156; 15'd5315: duty=145; 15'd5316: duty=140; 15'd5317: duty=141; 15'd5318: duty=129; 15'd5319: duty=127;
15'd5320: duty=129; 15'd5321: duty=131; 15'd5322: duty=132; 15'd5323: duty=127; 15'd5324: duty=129; 15'd5325: duty=120; 15'd5326: duty=131; 15'd5327: duty=131;
15'd5328: duty=121; 15'd5329: duty=120; 15'd5330: duty=118; 15'd5331: duty=110; 15'd5332: duty=118; 15'd5333: duty=115; 15'd5334: duty=107; 15'd5335: duty=115;
15'd5336: duty=115; 15'd5337: duty=109; 15'd5338: duty=104; 15'd5339: duty=96; 15'd5340: duty=105; 15'd5341: duty=122; 15'd5342: duty=121; 15'd5343: duty=118;
15'd5344: duty=120; 15'd5345: duty=134; 15'd5346: duty=136; 15'd5347: duty=128; 15'd5348: duty=130; 15'd5349: duty=134; 15'd5350: duty=133; 15'd5351: duty=135;
15'd5352: duty=137; 15'd5353: duty=135; 15'd5354: duty=136; 15'd5355: duty=140; 15'd5356: duty=144; 15'd5357: duty=138; 15'd5358: duty=139; 15'd5359: duty=146;
15'd5360: duty=153; 15'd5361: duty=143; 15'd5362: duty=144; 15'd5363: duty=143; 15'd5364: duty=138; 15'd5365: duty=149; 15'd5366: duty=151; 15'd5367: duty=149;
15'd5368: duty=145; 15'd5369: duty=146; 15'd5370: duty=147; 15'd5371: duty=145; 15'd5372: duty=133; 15'd5373: duty=140; 15'd5374: duty=144; 15'd5375: duty=139;
15'd5376: duty=133; 15'd5377: duty=134; 15'd5378: duty=138; 15'd5379: duty=139; 15'd5380: duty=136; 15'd5381: duty=122; 15'd5382: duty=118; 15'd5383: duty=125;
15'd5384: duty=125; 15'd5385: duty=108; 15'd5386: duty=103; 15'd5387: duty=101; 15'd5388: duty=101; 15'd5389: duty=98; 15'd5390: duty=98; 15'd5391: duty=103;
15'd5392: duty=109; 15'd5393: duty=108; 15'd5394: duty=105; 15'd5395: duty=104; 15'd5396: duty=105; 15'd5397: duty=107; 15'd5398: duty=108; 15'd5399: duty=105;
15'd5400: duty=96; 15'd5401: duty=98; 15'd5402: duty=102; 15'd5403: duty=105; 15'd5404: duty=111; 15'd5405: duty=113; 15'd5406: duty=112; 15'd5407: duty=119;
15'd5408: duty=124; 15'd5409: duty=129; 15'd5410: duty=131; 15'd5411: duty=134; 15'd5412: duty=140; 15'd5413: duty=150; 15'd5414: duty=151; 15'd5415: duty=159;
15'd5416: duty=165; 15'd5417: duty=162; 15'd5418: duty=160; 15'd5419: duty=159; 15'd5420: duty=165; 15'd5421: duty=167; 15'd5422: duty=167; 15'd5423: duty=161;
15'd5424: duty=162; 15'd5425: duty=168; 15'd5426: duty=171; 15'd5427: duty=167; 15'd5428: duty=166; 15'd5429: duty=165; 15'd5430: duty=169; 15'd5431: duty=167;
15'd5432: duty=165; 15'd5433: duty=162; 15'd5434: duty=160; 15'd5435: duty=162; 15'd5436: duty=157; 15'd5437: duty=150; 15'd5438: duty=149; 15'd5439: duty=153;
15'd5440: duty=145; 15'd5441: duty=137; 15'd5442: duty=137; 15'd5443: duty=133; 15'd5444: duty=129; 15'd5445: duty=131; 15'd5446: duty=125; 15'd5447: duty=116;
15'd5448: duty=116; 15'd5449: duty=120; 15'd5450: duty=122; 15'd5451: duty=121; 15'd5452: duty=116; 15'd5453: duty=112; 15'd5454: duty=111; 15'd5455: duty=107;
15'd5456: duty=102; 15'd5457: duty=90; 15'd5458: duty=90; 15'd5459: duty=81; 15'd5460: duty=73; 15'd5461: duty=72; 15'd5462: duty=76; 15'd5463: duty=75;
15'd5464: duty=69; 15'd5465: duty=78; 15'd5466: duty=87; 15'd5467: duty=99; 15'd5468: duty=104; 15'd5469: duty=108; 15'd5470: duty=111; 15'd5471: duty=111;
15'd5472: duty=115; 15'd5473: duty=122; 15'd5474: duty=118; 15'd5475: duty=120; 15'd5476: duty=128; 15'd5477: duty=132; 15'd5478: duty=127; 15'd5479: duty=135;
15'd5480: duty=132; 15'd5481: duty=140; 15'd5482: duty=150; 15'd5483: duty=140; 15'd5484: duty=142; 15'd5485: duty=149; 15'd5486: duty=156; 15'd5487: duty=163;
15'd5488: duty=170; 15'd5489: duty=155; 15'd5490: duty=153; 15'd5491: duty=163; 15'd5492: duty=159; 15'd5493: duty=169; 15'd5494: duty=167; 15'd5495: duty=166;
15'd5496: duty=157; 15'd5497: duty=152; 15'd5498: duty=151; 15'd5499: duty=146; 15'd5500: duty=145; 15'd5501: duty=156; 15'd5502: duty=150; 15'd5503: duty=122;
15'd5504: duty=133; 15'd5505: duty=146; 15'd5506: duty=133; 15'd5507: duty=127; 15'd5508: duty=131; 15'd5509: duty=103; 15'd5510: duty=105; 15'd5511: duty=113;
15'd5512: duty=117; 15'd5513: duty=125; 15'd5514: duty=123; 15'd5515: duty=137; 15'd5516: duty=145; 15'd5517: duty=130; 15'd5518: duty=127; 15'd5519: duty=144;
15'd5520: duty=127; 15'd5521: duty=119; 15'd5522: duty=125; 15'd5523: duty=113; 15'd5524: duty=121; 15'd5525: duty=128; 15'd5526: duty=112; 15'd5527: duty=116;
15'd5528: duty=119; 15'd5529: duty=126; 15'd5530: duty=142; 15'd5531: duty=145; 15'd5532: duty=151; 15'd5533: duty=150; 15'd5534: duty=148; 15'd5535: duty=145;
15'd5536: duty=139; 15'd5537: duty=145; 15'd5538: duty=150; 15'd5539: duty=136; 15'd5540: duty=136; 15'd5541: duty=145; 15'd5542: duty=136; 15'd5543: duty=156;
15'd5544: duty=152; 15'd5545: duty=155; 15'd5546: duty=147; 15'd5547: duty=139; 15'd5548: duty=135; 15'd5549: duty=114; 15'd5550: duty=121; 15'd5551: duty=126;
15'd5552: duty=120; 15'd5553: duty=120; 15'd5554: duty=115; 15'd5555: duty=114; 15'd5556: duty=117; 15'd5557: duty=102; 15'd5558: duty=112; 15'd5559: duty=105;
15'd5560: duty=103; 15'd5561: duty=110; 15'd5562: duty=115; 15'd5563: duty=105; 15'd5564: duty=96; 15'd5565: duty=105; 15'd5566: duty=112; 15'd5567: duty=103;
15'd5568: duty=98; 15'd5569: duty=99; 15'd5570: duty=79; 15'd5571: duty=90; 15'd5572: duty=93; 15'd5573: duty=88; 15'd5574: duty=94; 15'd5575: duty=93;
15'd5576: duty=104; 15'd5577: duty=101; 15'd5578: duty=97; 15'd5579: duty=100; 15'd5580: duty=105; 15'd5581: duty=121; 15'd5582: duty=123; 15'd5583: duty=107;
15'd5584: duty=119; 15'd5585: duty=130; 15'd5586: duty=137; 15'd5587: duty=145; 15'd5588: duty=149; 15'd5589: duty=168; 15'd5590: duty=177; 15'd5591: duty=182;
15'd5592: duty=180; 15'd5593: duty=176; 15'd5594: duty=176; 15'd5595: duty=184; 15'd5596: duty=179; 15'd5597: duty=176; 15'd5598: duty=180; 15'd5599: duty=179;
15'd5600: duty=182; 15'd5601: duty=185; 15'd5602: duty=177; 15'd5603: duty=188; 15'd5604: duty=188; 15'd5605: duty=177; 15'd5606: duty=177; 15'd5607: duty=177;
15'd5608: duty=175; 15'd5609: duty=168; 15'd5610: duty=162; 15'd5611: duty=165; 15'd5612: duty=168; 15'd5613: duty=154; 15'd5614: duty=153; 15'd5615: duty=159;
15'd5616: duty=147; 15'd5617: duty=133; 15'd5618: duty=141; 15'd5619: duty=136; 15'd5620: duty=123; 15'd5621: duty=121; 15'd5622: duty=110; 15'd5623: duty=107;
15'd5624: duty=102; 15'd5625: duty=93; 15'd5626: duty=93; 15'd5627: duty=90; 15'd5628: duty=91; 15'd5629: duty=91; 15'd5630: duty=85; 15'd5631: duty=76;
15'd5632: duty=79; 15'd5633: duty=87; 15'd5634: duty=88; 15'd5635: duty=84; 15'd5636: duty=79; 15'd5637: duty=84; 15'd5638: duty=82; 15'd5639: duty=84;
15'd5640: duty=85; 15'd5641: duty=79; 15'd5642: duty=81; 15'd5643: duty=87; 15'd5644: duty=90; 15'd5645: duty=85; 15'd5646: duty=93; 15'd5647: duty=102;
15'd5648: duty=104; 15'd5649: duty=114; 15'd5650: duty=116; 15'd5651: duty=120; 15'd5652: duty=128; 15'd5653: duty=132; 15'd5654: duty=136; 15'd5655: duty=140;
15'd5656: duty=135; 15'd5657: duty=135; 15'd5658: duty=144; 15'd5659: duty=139; 15'd5660: duty=139; 15'd5661: duty=146; 15'd5662: duty=141; 15'd5663: duty=141;
15'd5664: duty=144; 15'd5665: duty=149; 15'd5666: duty=164; 15'd5667: duty=166; 15'd5668: duty=167; 15'd5669: duty=171; 15'd5670: duty=174; 15'd5671: duty=174;
15'd5672: duty=170; 15'd5673: duty=165; 15'd5674: duty=162; 15'd5675: duty=163; 15'd5676: duty=161; 15'd5677: duty=162; 15'd5678: duty=156; 15'd5679: duty=152;
15'd5680: duty=154; 15'd5681: duty=151; 15'd5682: duty=142; 15'd5683: duty=139; 15'd5684: duty=145; 15'd5685: duty=151; 15'd5686: duty=146; 15'd5687: duty=143;
15'd5688: duty=134; 15'd5689: duty=132; 15'd5690: duty=129; 15'd5691: duty=129; 15'd5692: duty=125; 15'd5693: duty=111; 15'd5694: duty=122; 15'd5695: duty=125;
15'd5696: duty=113; 15'd5697: duty=114; 15'd5698: duty=113; 15'd5699: duty=113; 15'd5700: duty=114; 15'd5701: duty=111; 15'd5702: duty=118; 15'd5703: duty=121;
15'd5704: duty=121; 15'd5705: duty=127; 15'd5706: duty=133; 15'd5707: duty=128; 15'd5708: duty=127; 15'd5709: duty=128; 15'd5710: duty=132; 15'd5711: duty=131;
15'd5712: duty=140; 15'd5713: duty=139; 15'd5714: duty=137; 15'd5715: duty=140; 15'd5716: duty=138; 15'd5717: duty=139; 15'd5718: duty=145; 15'd5719: duty=147;
15'd5720: duty=143; 15'd5721: duty=142; 15'd5722: duty=143; 15'd5723: duty=144; 15'd5724: duty=143; 15'd5725: duty=145; 15'd5726: duty=142; 15'd5727: duty=141;
15'd5728: duty=140; 15'd5729: duty=144; 15'd5730: duty=137; 15'd5731: duty=134; 15'd5732: duty=131; 15'd5733: duty=126; 15'd5734: duty=122; 15'd5735: duty=121;
15'd5736: duty=121; 15'd5737: duty=124; 15'd5738: duty=116; 15'd5739: duty=119; 15'd5740: duty=118; 15'd5741: duty=110; 15'd5742: duty=116; 15'd5743: duty=122;
15'd5744: duty=128; 15'd5745: duty=118; 15'd5746: duty=112; 15'd5747: duty=116; 15'd5748: duty=115; 15'd5749: duty=111; 15'd5750: duty=109; 15'd5751: duty=95;
15'd5752: duty=97; 15'd5753: duty=98; 15'd5754: duty=97; 15'd5755: duty=93; 15'd5756: duty=98; 15'd5757: duty=93; 15'd5758: duty=94; 15'd5759: duty=99;
15'd5760: duty=95; 15'd5761: duty=103; 15'd5762: duty=110; 15'd5763: duty=112; 15'd5764: duty=118; 15'd5765: duty=121; 15'd5766: duty=120; 15'd5767: duty=128;
15'd5768: duty=133; 15'd5769: duty=136; 15'd5770: duty=139; 15'd5771: duty=145; 15'd5772: duty=144; 15'd5773: duty=153; 15'd5774: duty=147; 15'd5775: duty=148;
15'd5776: duty=151; 15'd5777: duty=154; 15'd5778: duty=154; 15'd5779: duty=149; 15'd5780: duty=149; 15'd5781: duty=151; 15'd5782: duty=154; 15'd5783: duty=145;
15'd5784: duty=154; 15'd5785: duty=165; 15'd5786: duty=162; 15'd5787: duty=161; 15'd5788: duty=160; 15'd5789: duty=161; 15'd5790: duty=157; 15'd5791: duty=157;
15'd5792: duty=157; 15'd5793: duty=152; 15'd5794: duty=156; 15'd5795: duty=153; 15'd5796: duty=153; 15'd5797: duty=155; 15'd5798: duty=153; 15'd5799: duty=150;
15'd5800: duty=137; 15'd5801: duty=132; 15'd5802: duty=131; 15'd5803: duty=129; 15'd5804: duty=135; 15'd5805: duty=139; 15'd5806: duty=133; 15'd5807: duty=126;
15'd5808: duty=118; 15'd5809: duty=121; 15'd5810: duty=127; 15'd5811: duty=121; 15'd5812: duty=119; 15'd5813: duty=113; 15'd5814: duty=119; 15'd5815: duty=117;
15'd5816: duty=116; 15'd5817: duty=118; 15'd5818: duty=117; 15'd5819: duty=121; 15'd5820: duty=117; 15'd5821: duty=118; 15'd5822: duty=117; 15'd5823: duty=119;
15'd5824: duty=125; 15'd5825: duty=129; 15'd5826: duty=134; 15'd5827: duty=124; 15'd5828: duty=115; 15'd5829: duty=121; 15'd5830: duty=122; 15'd5831: duty=112;
15'd5832: duty=116; 15'd5833: duty=120; 15'd5834: duty=114; 15'd5835: duty=119; 15'd5836: duty=124; 15'd5837: duty=133; 15'd5838: duty=134; 15'd5839: duty=140;
15'd5840: duty=145; 15'd5841: duty=152; 15'd5842: duty=153; 15'd5843: duty=149; 15'd5844: duty=136; 15'd5845: duty=136; 15'd5846: duty=136; 15'd5847: duty=132;
15'd5848: duty=131; 15'd5849: duty=125; 15'd5850: duty=130; 15'd5851: duty=133; 15'd5852: duty=130; 15'd5853: duty=124; 15'd5854: duty=134; 15'd5855: duty=139;
15'd5856: duty=136; 15'd5857: duty=141; 15'd5858: duty=144; 15'd5859: duty=143; 15'd5860: duty=130; 15'd5861: duty=111; 15'd5862: duty=115; 15'd5863: duty=105;
15'd5864: duty=89; 15'd5865: duty=93; 15'd5866: duty=90; 15'd5867: duty=81; 15'd5868: duty=78; 15'd5869: duty=82; 15'd5870: duty=95; 15'd5871: duty=101;
15'd5872: duty=107; 15'd5873: duty=116; 15'd5874: duty=123; 15'd5875: duty=122; 15'd5876: duty=122; 15'd5877: duty=131; 15'd5878: duty=127; 15'd5879: duty=116;
15'd5880: duty=109; 15'd5881: duty=121; 15'd5882: duty=113; 15'd5883: duty=122; 15'd5884: duty=124; 15'd5885: duty=124; 15'd5886: duty=145; 15'd5887: duty=134;
15'd5888: duty=150; 15'd5889: duty=160; 15'd5890: duty=156; 15'd5891: duty=162; 15'd5892: duty=167; 15'd5893: duty=174; 15'd5894: duty=173; 15'd5895: duty=175;
15'd5896: duty=182; 15'd5897: duty=176; 15'd5898: duty=172; 15'd5899: duty=180; 15'd5900: duty=170; 15'd5901: duty=176; 15'd5902: duty=171; 15'd5903: duty=172;
15'd5904: duty=181; 15'd5905: duty=169; 15'd5906: duty=161; 15'd5907: duty=154; 15'd5908: duty=157; 15'd5909: duty=149; 15'd5910: duty=144; 15'd5911: duty=138;
15'd5912: duty=134; 15'd5913: duty=136; 15'd5914: duty=128; 15'd5915: duty=132; 15'd5916: duty=141; 15'd5917: duty=127; 15'd5918: duty=128; 15'd5919: duty=130;
15'd5920: duty=124; 15'd5921: duty=119; 15'd5922: duty=118; 15'd5923: duty=130; 15'd5924: duty=122; 15'd5925: duty=121; 15'd5926: duty=117; 15'd5927: duty=98;
15'd5928: duty=95; 15'd5929: duty=95; 15'd5930: duty=98; 15'd5931: duty=98; 15'd5932: duty=99; 15'd5933: duty=107; 15'd5934: duty=110; 15'd5935: duty=114;
15'd5936: duty=113; 15'd5937: duty=107; 15'd5938: duty=108; 15'd5939: duty=112; 15'd5940: duty=102; 15'd5941: duty=102; 15'd5942: duty=98; 15'd5943: duty=92;
15'd5944: duty=92; 15'd5945: duty=93; 15'd5946: duty=92; 15'd5947: duty=99; 15'd5948: duty=117; 15'd5949: duty=124; 15'd5950: duty=131; 15'd5951: duty=141;
15'd5952: duty=143; 15'd5953: duty=148; 15'd5954: duty=148; 15'd5955: duty=144; 15'd5956: duty=151; 15'd5957: duty=145; 15'd5958: duty=138; 15'd5959: duty=142;
15'd5960: duty=137; 15'd5961: duty=129; 15'd5962: duty=137; 15'd5963: duty=138; 15'd5964: duty=136; 15'd5965: duty=139; 15'd5966: duty=153; 15'd5967: duty=150;
15'd5968: duty=145; 15'd5969: duty=154; 15'd5970: duty=148; 15'd5971: duty=149; 15'd5972: duty=149; 15'd5973: duty=150; 15'd5974: duty=140; 15'd5975: duty=135;
15'd5976: duty=138; 15'd5977: duty=134; 15'd5978: duty=125; 15'd5979: duty=120; 15'd5980: duty=119; 15'd5981: duty=125; 15'd5982: duty=124; 15'd5983: duty=116;
15'd5984: duty=120; 15'd5985: duty=122; 15'd5986: duty=122; 15'd5987: duty=122; 15'd5988: duty=121; 15'd5989: duty=120; 15'd5990: duty=118; 15'd5991: duty=120;
15'd5992: duty=127; 15'd5993: duty=125; 15'd5994: duty=124; 15'd5995: duty=128; 15'd5996: duty=130; 15'd5997: duty=134; 15'd5998: duty=129; 15'd5999: duty=130;
15'd6000: duty=133; 15'd6001: duty=133; 15'd6002: duty=142; 15'd6003: duty=142; 15'd6004: duty=139; 15'd6005: duty=153; 15'd6006: duty=159; 15'd6007: duty=163;
15'd6008: duty=164; 15'd6009: duty=154; 15'd6010: duty=159; 15'd6011: duty=167; 15'd6012: duty=160; 15'd6013: duty=153; 15'd6014: duty=156; 15'd6015: duty=143;
15'd6016: duty=136; 15'd6017: duty=136; 15'd6018: duty=130; 15'd6019: duty=131; 15'd6020: duty=138; 15'd6021: duty=137; 15'd6022: duty=137; 15'd6023: duty=146;
15'd6024: duty=155; 15'd6025: duty=160; 15'd6026: duty=152; 15'd6027: duty=151; 15'd6028: duty=153; 15'd6029: duty=146; 15'd6030: duty=135; 15'd6031: duty=131;
15'd6032: duty=129; 15'd6033: duty=122; 15'd6034: duty=109; 15'd6035: duty=104; 15'd6036: duty=96; 15'd6037: duty=93; 15'd6038: duty=98; 15'd6039: duty=95;
15'd6040: duty=96; 15'd6041: duty=102; 15'd6042: duty=98; 15'd6043: duty=101; 15'd6044: duty=105; 15'd6045: duty=100; 15'd6046: duty=93; 15'd6047: duty=98;
15'd6048: duty=101; 15'd6049: duty=101; 15'd6050: duty=96; 15'd6051: duty=92; 15'd6052: duty=96; 15'd6053: duty=100; 15'd6054: duty=98; 15'd6055: duty=92;
15'd6056: duty=95; 15'd6057: duty=101; 15'd6058: duty=106; 15'd6059: duty=106; 15'd6060: duty=111; 15'd6061: duty=112; 15'd6062: duty=128; 15'd6063: duty=128;
15'd6064: duty=134; 15'd6065: duty=133; 15'd6066: duty=135; 15'd6067: duty=138; 15'd6068: duty=145; 15'd6069: duty=152; 15'd6070: duty=154; 15'd6071: duty=157;
15'd6072: duty=160; 15'd6073: duty=158; 15'd6074: duty=158; 15'd6075: duty=169; 15'd6076: duty=167; 15'd6077: duty=171; 15'd6078: duty=177; 15'd6079: duty=180;
15'd6080: duty=174; 15'd6081: duty=176; 15'd6082: duty=169; 15'd6083: duty=169; 15'd6084: duty=160; 15'd6085: duty=159; 15'd6086: duty=160; 15'd6087: duty=159;
15'd6088: duty=155; 15'd6089: duty=153; 15'd6090: duty=160; 15'd6091: duty=157; 15'd6092: duty=149; 15'd6093: duty=150; 15'd6094: duty=151; 15'd6095: duty=147;
15'd6096: duty=144; 15'd6097: duty=136; 15'd6098: duty=128; 15'd6099: duty=127; 15'd6100: duty=130; 15'd6101: duty=124; 15'd6102: duty=116; 15'd6103: duty=110;
15'd6104: duty=121; 15'd6105: duty=118; 15'd6106: duty=117; 15'd6107: duty=109; 15'd6108: duty=103; 15'd6109: duty=112; 15'd6110: duty=109; 15'd6111: duty=98;
15'd6112: duty=105; 15'd6113: duty=103; 15'd6114: duty=104; 15'd6115: duty=104; 15'd6116: duty=104; 15'd6117: duty=106; 15'd6118: duty=104; 15'd6119: duty=107;
15'd6120: duty=107; 15'd6121: duty=104; 15'd6122: duty=102; 15'd6123: duty=116; 15'd6124: duty=114; 15'd6125: duty=115; 15'd6126: duty=120; 15'd6127: duty=121;
15'd6128: duty=121; 15'd6129: duty=121; 15'd6130: duty=119; 15'd6131: duty=124; 15'd6132: duty=127; 15'd6133: duty=130; 15'd6134: duty=131; 15'd6135: duty=134;
15'd6136: duty=128; 15'd6137: duty=128; 15'd6138: duty=131; 15'd6139: duty=136; 15'd6140: duty=134; 15'd6141: duty=130; 15'd6142: duty=137; 15'd6143: duty=136;
15'd6144: duty=143; 15'd6145: duty=142; 15'd6146: duty=140; 15'd6147: duty=137; 15'd6148: duty=131; 15'd6149: duty=137; 15'd6150: duty=140; 15'd6151: duty=135;
15'd6152: duty=140; 15'd6153: duty=137; 15'd6154: duty=139; 15'd6155: duty=137; 15'd6156: duty=134; 15'd6157: duty=134; 15'd6158: duty=128; 15'd6159: duty=126;
15'd6160: duty=128; 15'd6161: duty=131; 15'd6162: duty=127; 15'd6163: duty=131; 15'd6164: duty=136; 15'd6165: duty=129; 15'd6166: duty=129; 15'd6167: duty=130;
15'd6168: duty=125; 15'd6169: duty=125; 15'd6170: duty=123; 15'd6171: duty=124; 15'd6172: duty=125; 15'd6173: duty=124; 15'd6174: duty=125; 15'd6175: duty=133;
15'd6176: duty=129; 15'd6177: duty=129; 15'd6178: duty=132; 15'd6179: duty=135; 15'd6180: duty=140; 15'd6181: duty=131; 15'd6182: duty=136; 15'd6183: duty=139;
15'd6184: duty=142; 15'd6185: duty=151; 15'd6186: duty=156; 15'd6187: duty=148; 15'd6188: duty=148; 15'd6189: duty=157; 15'd6190: duty=153; 15'd6191: duty=151;
15'd6192: duty=157; 15'd6193: duty=157; 15'd6194: duty=154; 15'd6195: duty=157; 15'd6196: duty=156; 15'd6197: duty=152; 15'd6198: duty=153; 15'd6199: duty=152;
15'd6200: duty=150; 15'd6201: duty=150; 15'd6202: duty=139; 15'd6203: duty=142; 15'd6204: duty=145; 15'd6205: duty=139; 15'd6206: duty=131; 15'd6207: duty=127;
15'd6208: duty=127; 15'd6209: duty=123; 15'd6210: duty=124; 15'd6211: duty=116; 15'd6212: duty=111; 15'd6213: duty=116; 15'd6214: duty=113; 15'd6215: duty=115;
15'd6216: duty=122; 15'd6217: duty=110; 15'd6218: duty=112; 15'd6219: duty=119; 15'd6220: duty=106; 15'd6221: duty=109; 15'd6222: duty=112; 15'd6223: duty=101;
15'd6224: duty=100; 15'd6225: duty=100; 15'd6226: duty=93; 15'd6227: duty=87; 15'd6228: duty=86; 15'd6229: duty=90; 15'd6230: duty=87; 15'd6231: duty=90;
15'd6232: duty=92; 15'd6233: duty=100; 15'd6234: duty=101; 15'd6235: duty=99; 15'd6236: duty=109; 15'd6237: duty=107; 15'd6238: duty=104; 15'd6239: duty=105;
15'd6240: duty=113; 15'd6241: duty=112; 15'd6242: duty=118; 15'd6243: duty=123; 15'd6244: duty=121; 15'd6245: duty=126; 15'd6246: duty=130; 15'd6247: duty=131;
15'd6248: duty=134; 15'd6249: duty=138; 15'd6250: duty=143; 15'd6251: duty=149; 15'd6252: duty=154; 15'd6253: duty=163; 15'd6254: duty=164; 15'd6255: duty=169;
15'd6256: duty=168; 15'd6257: duty=168; 15'd6258: duty=167; 15'd6259: duty=166; 15'd6260: duty=171; 15'd6261: duty=176; 15'd6262: duty=168; 15'd6263: duty=167;
15'd6264: duty=171; 15'd6265: duty=167; 15'd6266: duty=167; 15'd6267: duty=164; 15'd6268: duty=164; 15'd6269: duty=166; 15'd6270: duty=164; 15'd6271: duty=160;
15'd6272: duty=157; 15'd6273: duty=156; 15'd6274: duty=148; 15'd6275: duty=143; 15'd6276: duty=137; 15'd6277: duty=135; 15'd6278: duty=136; 15'd6279: duty=129;
15'd6280: duty=129; 15'd6281: duty=131; 15'd6282: duty=127; 15'd6283: duty=129; 15'd6284: duty=128; 15'd6285: duty=127; 15'd6286: duty=128; 15'd6287: duty=122;
15'd6288: duty=116; 15'd6289: duty=113; 15'd6290: duty=113; 15'd6291: duty=110; 15'd6292: duty=109; 15'd6293: duty=104; 15'd6294: duty=106; 15'd6295: duty=107;
15'd6296: duty=104; 15'd6297: duty=112; 15'd6298: duty=110; 15'd6299: duty=105; 15'd6300: duty=111; 15'd6301: duty=112; 15'd6302: duty=112; 15'd6303: duty=118;
15'd6304: duty=120; 15'd6305: duty=121; 15'd6306: duty=126; 15'd6307: duty=132; 15'd6308: duty=131; 15'd6309: duty=130; 15'd6310: duty=131; 15'd6311: duty=139;
15'd6312: duty=141; 15'd6313: duty=139; 15'd6314: duty=137; 15'd6315: duty=136; 15'd6316: duty=129; 15'd6317: duty=119; 15'd6318: duty=119; 15'd6319: duty=122;
15'd6320: duty=124; 15'd6321: duty=121; 15'd6322: duty=119; 15'd6323: duty=115; 15'd6324: duty=116; 15'd6325: duty=121; 15'd6326: duty=125; 15'd6327: duty=128;
15'd6328: duty=125; 15'd6329: duty=129; 15'd6330: duty=135; 15'd6331: duty=133; 15'd6332: duty=135; 15'd6333: duty=132; 15'd6334: duty=137; 15'd6335: duty=136;
15'd6336: duty=128; 15'd6337: duty=131; 15'd6338: duty=121; 15'd6339: duty=127; 15'd6340: duty=129; 15'd6341: duty=119; 15'd6342: duty=118; 15'd6343: duty=118;
15'd6344: duty=115; 15'd6345: duty=116; 15'd6346: duty=121; 15'd6347: duty=128; 15'd6348: duty=131; 15'd6349: duty=128; 15'd6350: duty=134; 15'd6351: duty=139;
15'd6352: duty=136; 15'd6353: duty=131; 15'd6354: duty=136; 15'd6355: duty=136; 15'd6356: duty=130; 15'd6357: duty=128; 15'd6358: duty=124; 15'd6359: duty=124;
15'd6360: duty=131; 15'd6361: duty=127; 15'd6362: duty=125; 15'd6363: duty=131; 15'd6364: duty=134; 15'd6365: duty=140; 15'd6366: duty=136; 15'd6367: duty=141;
15'd6368: duty=150; 15'd6369: duty=150; 15'd6370: duty=151; 15'd6371: duty=156; 15'd6372: duty=159; 15'd6373: duty=161; 15'd6374: duty=159; 15'd6375: duty=159;
15'd6376: duty=154; 15'd6377: duty=148; 15'd6378: duty=156; 15'd6379: duty=156; 15'd6380: duty=151; 15'd6381: duty=145; 15'd6382: duty=141; 15'd6383: duty=143;
15'd6384: duty=148; 15'd6385: duty=143; 15'd6386: duty=142; 15'd6387: duty=142; 15'd6388: duty=137; 15'd6389: duty=140; 15'd6390: duty=137; 15'd6391: duty=131;
15'd6392: duty=129; 15'd6393: duty=130; 15'd6394: duty=122; 15'd6395: duty=121; 15'd6396: duty=118; 15'd6397: duty=113; 15'd6398: duty=121; 15'd6399: duty=125;
15'd6400: duty=122; 15'd6401: duty=122; 15'd6402: duty=125; 15'd6403: duty=127; 15'd6404: duty=128; 15'd6405: duty=123; 15'd6406: duty=119; 15'd6407: duty=121;
15'd6408: duty=113; 15'd6409: duty=109; 15'd6410: duty=109; 15'd6411: duty=107; 15'd6412: duty=105; 15'd6413: duty=106; 15'd6414: duty=108; 15'd6415: duty=104;
15'd6416: duty=107; 15'd6417: duty=113; 15'd6418: duty=112; 15'd6419: duty=109; 15'd6420: duty=114; 15'd6421: duty=112; 15'd6422: duty=118; 15'd6423: duty=121;
15'd6424: duty=118; 15'd6425: duty=121; 15'd6426: duty=121; 15'd6427: duty=128; 15'd6428: duty=130; 15'd6429: duty=129; 15'd6430: duty=125; 15'd6431: duty=125;
15'd6432: duty=130; 15'd6433: duty=129; 15'd6434: duty=131; 15'd6435: duty=131; 15'd6436: duty=134; 15'd6437: duty=137; 15'd6438: duty=139; 15'd6439: duty=139;
15'd6440: duty=140; 15'd6441: duty=143; 15'd6442: duty=146; 15'd6443: duty=143; 15'd6444: duty=139; 15'd6445: duty=142; 15'd6446: duty=147; 15'd6447: duty=143;
15'd6448: duty=143; 15'd6449: duty=144; 15'd6450: duty=144; 15'd6451: duty=139; 15'd6452: duty=134; 15'd6453: duty=137; 15'd6454: duty=136; 15'd6455: duty=136;
15'd6456: duty=139; 15'd6457: duty=140; 15'd6458: duty=140; 15'd6459: duty=140; 15'd6460: duty=141; 15'd6461: duty=142; 15'd6462: duty=140; 15'd6463: duty=137;
15'd6464: duty=134; 15'd6465: duty=127; 15'd6466: duty=128; 15'd6467: duty=130; 15'd6468: duty=118; 15'd6469: duty=125; 15'd6470: duty=124; 15'd6471: duty=132;
15'd6472: duty=133; 15'd6473: duty=129; 15'd6474: duty=133; 15'd6475: duty=134; 15'd6476: duty=131; 15'd6477: duty=124; 15'd6478: duty=127; 15'd6479: duty=131;
15'd6480: duty=128; 15'd6481: duty=126; 15'd6482: duty=126; 15'd6483: duty=121; 15'd6484: duty=124; 15'd6485: duty=136; 15'd6486: duty=142; 15'd6487: duty=142;
15'd6488: duty=140; 15'd6489: duty=142; 15'd6490: duty=143; 15'd6491: duty=143; 15'd6492: duty=135; 15'd6493: duty=136; 15'd6494: duty=146; 15'd6495: duty=145;
15'd6496: duty=148; 15'd6497: duty=142; 15'd6498: duty=147; 15'd6499: duty=144; 15'd6500: duty=139; 15'd6501: duty=134; 15'd6502: duty=133; 15'd6503: duty=137;
15'd6504: duty=139; 15'd6505: duty=128; 15'd6506: duty=127; 15'd6507: duty=125; 15'd6508: duty=124; 15'd6509: duty=127; 15'd6510: duty=124; 15'd6511: duty=139;
15'd6512: duty=131; 15'd6513: duty=127; 15'd6514: duty=127; 15'd6515: duty=127; 15'd6516: duty=115; 15'd6517: duty=98; 15'd6518: duty=104; 15'd6519: duty=109;
15'd6520: duty=98; 15'd6521: duty=91; 15'd6522: duty=87; 15'd6523: duty=101; 15'd6524: duty=109; 15'd6525: duty=99; 15'd6526: duty=107; 15'd6527: duty=105;
15'd6528: duty=104; 15'd6529: duty=112; 15'd6530: duty=102; 15'd6531: duty=101; 15'd6532: duty=101; 15'd6533: duty=99; 15'd6534: duty=104; 15'd6535: duty=106;
15'd6536: duty=108; 15'd6537: duty=109; 15'd6538: duty=119; 15'd6539: duty=124; 15'd6540: duty=130; 15'd6541: duty=144; 15'd6542: duty=142; 15'd6543: duty=147;
15'd6544: duty=151; 15'd6545: duty=139; 15'd6546: duty=131; 15'd6547: duty=140; 15'd6548: duty=150; 15'd6549: duty=153; 15'd6550: duty=160; 15'd6551: duty=152;
15'd6552: duty=151; 15'd6553: duty=165; 15'd6554: duty=171; 15'd6555: duty=174; 15'd6556: duty=177; 15'd6557: duty=184; 15'd6558: duty=182; 15'd6559: duty=179;
15'd6560: duty=175; 15'd6561: duty=174; 15'd6562: duty=182; 15'd6563: duty=176; 15'd6564: duty=167; 15'd6565: duty=166; 15'd6566: duty=158; 15'd6567: duty=157;
15'd6568: duty=165; 15'd6569: duty=155; 15'd6570: duty=145; 15'd6571: duty=137; 15'd6572: duty=138; 15'd6573: duty=137; 15'd6574: duty=131; 15'd6575: duty=135;
15'd6576: duty=127; 15'd6577: duty=121; 15'd6578: duty=127; 15'd6579: duty=120; 15'd6580: duty=116; 15'd6581: duty=110; 15'd6582: duty=109; 15'd6583: duty=114;
15'd6584: duty=106; 15'd6585: duty=96; 15'd6586: duty=92; 15'd6587: duty=87; 15'd6588: duty=89; 15'd6589: duty=90; 15'd6590: duty=87; 15'd6591: duty=88;
15'd6592: duty=93; 15'd6593: duty=101; 15'd6594: duty=89; 15'd6595: duty=93; 15'd6596: duty=92; 15'd6597: duty=88; 15'd6598: duty=95; 15'd6599: duty=91;
15'd6600: duty=86; 15'd6601: duty=88; 15'd6602: duty=84; 15'd6603: duty=94; 15'd6604: duty=103; 15'd6605: duty=102; 15'd6606: duty=110; 15'd6607: duty=124;
15'd6608: duty=140; 15'd6609: duty=140; 15'd6610: duty=151; 15'd6611: duty=159; 15'd6612: duty=153; 15'd6613: duty=154; 15'd6614: duty=154; 15'd6615: duty=153;
15'd6616: duty=159; 15'd6617: duty=157; 15'd6618: duty=157; 15'd6619: duty=157; 15'd6620: duty=159; 15'd6621: duty=165; 15'd6622: duty=164; 15'd6623: duty=160;
15'd6624: duty=166; 15'd6625: duty=167; 15'd6626: duty=165; 15'd6627: duty=162; 15'd6628: duty=171; 15'd6629: duty=166; 15'd6630: duty=164; 15'd6631: duty=162;
15'd6632: duty=162; 15'd6633: duty=162; 15'd6634: duty=154; 15'd6635: duty=148; 15'd6636: duty=142; 15'd6637: duty=137; 15'd6638: duty=128; 15'd6639: duty=124;
15'd6640: duty=119; 15'd6641: duty=116; 15'd6642: duty=111; 15'd6643: duty=116; 15'd6644: duty=114; 15'd6645: duty=113; 15'd6646: duty=108; 15'd6647: duty=113;
15'd6648: duty=121; 15'd6649: duty=123; 15'd6650: duty=121; 15'd6651: duty=121; 15'd6652: duty=112; 15'd6653: duty=102; 15'd6654: duty=108; 15'd6655: duty=107;
15'd6656: duty=105; 15'd6657: duty=96; 15'd6658: duty=95; 15'd6659: duty=98; 15'd6660: duty=99; 15'd6661: duty=99; 15'd6662: duty=102; 15'd6663: duty=106;
15'd6664: duty=119; 15'd6665: duty=125; 15'd6666: duty=125; 15'd6667: duty=128; 15'd6668: duty=134; 15'd6669: duty=139; 15'd6670: duty=143; 15'd6671: duty=150;
15'd6672: duty=145; 15'd6673: duty=142; 15'd6674: duty=148; 15'd6675: duty=148; 15'd6676: duty=149; 15'd6677: duty=147; 15'd6678: duty=146; 15'd6679: duty=142;
15'd6680: duty=148; 15'd6681: duty=157; 15'd6682: duty=156; 15'd6683: duty=159; 15'd6684: duty=160; 15'd6685: duty=162; 15'd6686: duty=158; 15'd6687: duty=162;
15'd6688: duty=163; 15'd6689: duty=157; 15'd6690: duty=148; 15'd6691: duty=144; 15'd6692: duty=137; 15'd6693: duty=133; 15'd6694: duty=137; 15'd6695: duty=134;
15'd6696: duty=127; 15'd6697: duty=127; 15'd6698: duty=129; 15'd6699: duty=130; 15'd6700: duty=132; 15'd6701: duty=127; 15'd6702: duty=125; 15'd6703: duty=127;
15'd6704: duty=121; 15'd6705: duty=115; 15'd6706: duty=112; 15'd6707: duty=101; 15'd6708: duty=93; 15'd6709: duty=92; 15'd6710: duty=101; 15'd6711: duty=95;
15'd6712: duty=93; 15'd6713: duty=105; 15'd6714: duty=108; 15'd6715: duty=108; 15'd6716: duty=104; 15'd6717: duty=110; 15'd6718: duty=117; 15'd6719: duty=109;
15'd6720: duty=113; 15'd6721: duty=110; 15'd6722: duty=104; 15'd6723: duty=109; 15'd6724: duty=113; 15'd6725: duty=116; 15'd6726: duty=116; 15'd6727: duty=122;
15'd6728: duty=127; 15'd6729: duty=137; 15'd6730: duty=148; 15'd6731: duty=146; 15'd6732: duty=146; 15'd6733: duty=148; 15'd6734: duty=145; 15'd6735: duty=146;
15'd6736: duty=142; 15'd6737: duty=145; 15'd6738: duty=145; 15'd6739: duty=148; 15'd6740: duty=156; 15'd6741: duty=153; 15'd6742: duty=157; 15'd6743: duty=164;
15'd6744: duty=170; 15'd6745: duty=168; 15'd6746: duty=166; 15'd6747: duty=167; 15'd6748: duty=169; 15'd6749: duty=167; 15'd6750: duty=166; 15'd6751: duty=160;
15'd6752: duty=151; 15'd6753: duty=153; 15'd6754: duty=154; 15'd6755: duty=148; 15'd6756: duty=138; 15'd6757: duty=141; 15'd6758: duty=139; 15'd6759: duty=136;
15'd6760: duty=132; 15'd6761: duty=119; 15'd6762: duty=118; 15'd6763: duty=123; 15'd6764: duty=121; 15'd6765: duty=115; 15'd6766: duty=114; 15'd6767: duty=127;
15'd6768: duty=124; 15'd6769: duty=118; 15'd6770: duty=110; 15'd6771: duty=106; 15'd6772: duty=104; 15'd6773: duty=101; 15'd6774: duty=94; 15'd6775: duty=82;
15'd6776: duty=87; 15'd6777: duty=90; 15'd6778: duty=93; 15'd6779: duty=84; 15'd6780: duty=84; 15'd6781: duty=89; 15'd6782: duty=93; 15'd6783: duty=99;
15'd6784: duty=99; 15'd6785: duty=101; 15'd6786: duty=104; 15'd6787: duty=113; 15'd6788: duty=118; 15'd6789: duty=116; 15'd6790: duty=122; 15'd6791: duty=119;
15'd6792: duty=128; 15'd6793: duty=131; 15'd6794: duty=134; 15'd6795: duty=137; 15'd6796: duty=138; 15'd6797: duty=142; 15'd6798: duty=142; 15'd6799: duty=145;
15'd6800: duty=147; 15'd6801: duty=154; 15'd6802: duty=159; 15'd6803: duty=162; 15'd6804: duty=153; 15'd6805: duty=158; 15'd6806: duty=164; 15'd6807: duty=168;
15'd6808: duty=177; 15'd6809: duty=169; 15'd6810: duty=167; 15'd6811: duty=174; 15'd6812: duty=170; 15'd6813: duty=167; 15'd6814: duty=165; 15'd6815: duty=165;
15'd6816: duty=161; 15'd6817: duty=162; 15'd6818: duty=160; 15'd6819: duty=154; 15'd6820: duty=151; 15'd6821: duty=150; 15'd6822: duty=152; 15'd6823: duty=148;
15'd6824: duty=147; 15'd6825: duty=142; 15'd6826: duty=142; 15'd6827: duty=142; 15'd6828: duty=132; 15'd6829: duty=128; 15'd6830: duty=122; 15'd6831: duty=118;
15'd6832: duty=115; 15'd6833: duty=106; 15'd6834: duty=109; 15'd6835: duty=110; 15'd6836: duty=107; 15'd6837: duty=107; 15'd6838: duty=107; 15'd6839: duty=96;
15'd6840: duty=99; 15'd6841: duty=102; 15'd6842: duty=98; 15'd6843: duty=93; 15'd6844: duty=87; 15'd6845: duty=87; 15'd6846: duty=87; 15'd6847: duty=89;
15'd6848: duty=85; 15'd6849: duty=90; 15'd6850: duty=96; 15'd6851: duty=104; 15'd6852: duty=107; 15'd6853: duty=105; 15'd6854: duty=112; 15'd6855: duty=118;
15'd6856: duty=122; 15'd6857: duty=125; 15'd6858: duty=123; 15'd6859: duty=121; 15'd6860: duty=127; 15'd6861: duty=131; 15'd6862: duty=134; 15'd6863: duty=139;
15'd6864: duty=142; 15'd6865: duty=145; 15'd6866: duty=153; 15'd6867: duty=154; 15'd6868: duty=151; 15'd6869: duty=154; 15'd6870: duty=162; 15'd6871: duty=165;
15'd6872: duty=163; 15'd6873: duty=159; 15'd6874: duty=156; 15'd6875: duty=156; 15'd6876: duty=156; 15'd6877: duty=156; 15'd6878: duty=145; 15'd6879: duty=145;
15'd6880: duty=144; 15'd6881: duty=142; 15'd6882: duty=141; 15'd6883: duty=142; 15'd6884: duty=137; 15'd6885: duty=136; 15'd6886: duty=140; 15'd6887: duty=145;
15'd6888: duty=139; 15'd6889: duty=139; 15'd6890: duty=146; 15'd6891: duty=142; 15'd6892: duty=142; 15'd6893: duty=143; 15'd6894: duty=139; 15'd6895: duty=137;
15'd6896: duty=142; 15'd6897: duty=136; 15'd6898: duty=131; 15'd6899: duty=131; 15'd6900: duty=126; 15'd6901: duty=119; 15'd6902: duty=119; 15'd6903: duty=118;
15'd6904: duty=118; 15'd6905: duty=115; 15'd6906: duty=115; 15'd6907: duty=120; 15'd6908: duty=118; 15'd6909: duty=115; 15'd6910: duty=116; 15'd6911: duty=110;
15'd6912: duty=107; 15'd6913: duty=112; 15'd6914: duty=113; 15'd6915: duty=110; 15'd6916: duty=111; 15'd6917: duty=107; 15'd6918: duty=114; 15'd6919: duty=119;
15'd6920: duty=115; 15'd6921: duty=120; 15'd6922: duty=119; 15'd6923: duty=123; 15'd6924: duty=124; 15'd6925: duty=127; 15'd6926: duty=127; 15'd6927: duty=128;
15'd6928: duty=125; 15'd6929: duty=127; 15'd6930: duty=128; 15'd6931: duty=125; 15'd6932: duty=128; 15'd6933: duty=136; 15'd6934: duty=137; 15'd6935: duty=133;
15'd6936: duty=146; 15'd6937: duty=139; 15'd6938: duty=143; 15'd6939: duty=153; 15'd6940: duty=150; 15'd6941: duty=153; 15'd6942: duty=147; 15'd6943: duty=147;
15'd6944: duty=152; 15'd6945: duty=147; 15'd6946: duty=147; 15'd6947: duty=145; 15'd6948: duty=143; 15'd6949: duty=142; 15'd6950: duty=143; 15'd6951: duty=137;
15'd6952: duty=134; 15'd6953: duty=136; 15'd6954: duty=133; 15'd6955: duty=137; 15'd6956: duty=134; 15'd6957: duty=136; 15'd6958: duty=139; 15'd6959: duty=142;
15'd6960: duty=143; 15'd6961: duty=145; 15'd6962: duty=139; 15'd6963: duty=140; 15'd6964: duty=140; 15'd6965: duty=137; 15'd6966: duty=139; 15'd6967: duty=131;
15'd6968: duty=129; 15'd6969: duty=127; 15'd6970: duty=122; 15'd6971: duty=119; 15'd6972: duty=119; 15'd6973: duty=119; 15'd6974: duty=118; 15'd6975: duty=124;
15'd6976: duty=122; 15'd6977: duty=120; 15'd6978: duty=121; 15'd6979: duty=116; 15'd6980: duty=121; 15'd6981: duty=121; 15'd6982: duty=119; 15'd6983: duty=117;
15'd6984: duty=125; 15'd6985: duty=126; 15'd6986: duty=122; 15'd6987: duty=127; 15'd6988: duty=125; 15'd6989: duty=124; 15'd6990: duty=122; 15'd6991: duty=124;
15'd6992: duty=122; 15'd6993: duty=121; 15'd6994: duty=122; 15'd6995: duty=124; 15'd6996: duty=120; 15'd6997: duty=118; 15'd6998: duty=118; 15'd6999: duty=118;
15'd7000: duty=118; 15'd7001: duty=123; 15'd7002: duty=124; 15'd7003: duty=128; 15'd7004: duty=133; 15'd7005: duty=127; 15'd7006: duty=131; 15'd7007: duty=136;
15'd7008: duty=137; 15'd7009: duty=136; 15'd7010: duty=134; 15'd7011: duty=134; 15'd7012: duty=136; 15'd7013: duty=139; 15'd7014: duty=143; 15'd7015: duty=142;
15'd7016: duty=137; 15'd7017: duty=131; 15'd7018: duty=134; 15'd7019: duty=131; 15'd7020: duty=134; 15'd7021: duty=136; 15'd7022: duty=130; 15'd7023: duty=131;
15'd7024: duty=133; 15'd7025: duty=134; 15'd7026: duty=133; 15'd7027: duty=131; 15'd7028: duty=136; 15'd7029: duty=137; 15'd7030: duty=142; 15'd7031: duty=150;
15'd7032: duty=148; 15'd7033: duty=148; 15'd7034: duty=142; 15'd7035: duty=139; 15'd7036: duty=137; 15'd7037: duty=136; 15'd7038: duty=129; 15'd7039: duty=130;
15'd7040: duty=136; 15'd7041: duty=137; 15'd7042: duty=143; 15'd7043: duty=142; 15'd7044: duty=139; 15'd7045: duty=142; 15'd7046: duty=148; 15'd7047: duty=144;
15'd7048: duty=138; 15'd7049: duty=139; 15'd7050: duty=141; 15'd7051: duty=136; 15'd7052: duty=131; 15'd7053: duty=132; 15'd7054: duty=129; 15'd7055: duty=127;
15'd7056: duty=132; 15'd7057: duty=130; 15'd7058: duty=127; 15'd7059: duty=124; 15'd7060: duty=127; 15'd7061: duty=126; 15'd7062: duty=122; 15'd7063: duty=124;
15'd7064: duty=122; 15'd7065: duty=121; 15'd7066: duty=117; 15'd7067: duty=115; 15'd7068: duty=115; 15'd7069: duty=117; 15'd7070: duty=122; 15'd7071: duty=122;
15'd7072: duty=116; 15'd7073: duty=122; 15'd7074: duty=128; 15'd7075: duty=125; 15'd7076: duty=122; 15'd7077: duty=118; 15'd7078: duty=113; 15'd7079: duty=115;
15'd7080: duty=116; 15'd7081: duty=116; 15'd7082: duty=118; 15'd7083: duty=122; 15'd7084: duty=125; 15'd7085: duty=125; 15'd7086: duty=125; 15'd7087: duty=121;
15'd7088: duty=124; 15'd7089: duty=121; 15'd7090: duty=122; 15'd7091: duty=119; 15'd7092: duty=110; 15'd7093: duty=111; 15'd7094: duty=109; 15'd7095: duty=107;
15'd7096: duty=107; 15'd7097: duty=115; 15'd7098: duty=121; 15'd7099: duty=126; 15'd7100: duty=133; 15'd7101: duty=137; 15'd7102: duty=137; 15'd7103: duty=140;
15'd7104: duty=143; 15'd7105: duty=145; 15'd7106: duty=148; 15'd7107: duty=156; 15'd7108: duty=157; 15'd7109: duty=161; 15'd7110: duty=159; 15'd7111: duty=153;
15'd7112: duty=151; 15'd7113: duty=150; 15'd7114: duty=154; 15'd7115: duty=148; 15'd7116: duty=154; 15'd7117: duty=150; 15'd7118: duty=151; 15'd7119: duty=156;
15'd7120: duty=152; 15'd7121: duty=154; 15'd7122: duty=157; 15'd7123: duty=158; 15'd7124: duty=155; 15'd7125: duty=154; 15'd7126: duty=145; 15'd7127: duty=138;
15'd7128: duty=137; 15'd7129: duty=133; 15'd7130: duty=141; 15'd7131: duty=134; 15'd7132: duty=125; 15'd7133: duty=121; 15'd7134: duty=119; 15'd7135: duty=128;
15'd7136: duty=119; 15'd7137: duty=121; 15'd7138: duty=128; 15'd7139: duty=124; 15'd7140: duty=119; 15'd7141: duty=120; 15'd7142: duty=114; 15'd7143: duty=109;
15'd7144: duty=114; 15'd7145: duty=115; 15'd7146: duty=111; 15'd7147: duty=112; 15'd7148: duty=108; 15'd7149: duty=107; 15'd7150: duty=105; 15'd7151: duty=101;
15'd7152: duty=102; 15'd7153: duty=98; 15'd7154: duty=99; 15'd7155: duty=112; 15'd7156: duty=121; 15'd7157: duty=122; 15'd7158: duty=127; 15'd7159: duty=134;
15'd7160: duty=135; 15'd7161: duty=137; 15'd7162: duty=136; 15'd7163: duty=142; 15'd7164: duty=142; 15'd7165: duty=140; 15'd7166: duty=142; 15'd7167: duty=128;
15'd7168: duty=128; 15'd7169: duty=121; 15'd7170: duty=119; 15'd7171: duty=126; 15'd7172: duty=129; 15'd7173: duty=139; 15'd7174: duty=146; 15'd7175: duty=143;
15'd7176: duty=151; 15'd7177: duty=151; 15'd7178: duty=157; 15'd7179: duty=165; 15'd7180: duty=164; 15'd7181: duty=157; 15'd7182: duty=148; 15'd7183: duty=143;
15'd7184: duty=144; 15'd7185: duty=139; 15'd7186: duty=130; 15'd7187: duty=134; 15'd7188: duty=131; 15'd7189: duty=133; 15'd7190: duty=131; 15'd7191: duty=131;
15'd7192: duty=134; 15'd7193: duty=137; 15'd7194: duty=131; 15'd7195: duty=132; 15'd7196: duty=133; 15'd7197: duty=131; 15'd7198: duty=126; 15'd7199: duty=119;
15'd7200: duty=115; 15'd7201: duty=111; 15'd7202: duty=109; 15'd7203: duty=117; 15'd7204: duty=116; 15'd7205: duty=114; 15'd7206: duty=117; 15'd7207: duty=113;
15'd7208: duty=112; 15'd7209: duty=113; 15'd7210: duty=110; 15'd7211: duty=104; 15'd7212: duty=115; 15'd7213: duty=111; 15'd7214: duty=109; 15'd7215: duty=117;
15'd7216: duty=119; 15'd7217: duty=114; 15'd7218: duty=112; 15'd7219: duty=116; 15'd7220: duty=118; 15'd7221: duty=117; 15'd7222: duty=124; 15'd7223: duty=124;
15'd7224: duty=118; 15'd7225: duty=122; 15'd7226: duty=130; 15'd7227: duty=134; 15'd7228: duty=135; 15'd7229: duty=149; 15'd7230: duty=155; 15'd7231: duty=158;
15'd7232: duty=164; 15'd7233: duty=171; 15'd7234: duty=170; 15'd7235: duty=171; 15'd7236: duty=176; 15'd7237: duty=163; 15'd7238: duty=158; 15'd7239: duty=162;
15'd7240: duty=153; 15'd7241: duty=146; 15'd7242: duty=145; 15'd7243: duty=149; 15'd7244: duty=150; 15'd7245: duty=152; 15'd7246: duty=150; 15'd7247: duty=155;
15'd7248: duty=161; 15'd7249: duty=157; 15'd7250: duty=158; 15'd7251: duty=152; 15'd7252: duty=156; 15'd7253: duty=155; 15'd7254: duty=151; 15'd7255: duty=145;
15'd7256: duty=134; 15'd7257: duty=129; 15'd7258: duty=127; 15'd7259: duty=122; 15'd7260: duty=115; 15'd7261: duty=108; 15'd7262: duty=107; 15'd7263: duty=108;
15'd7264: duty=104; 15'd7265: duty=99; 15'd7266: duty=100; 15'd7267: duty=102; 15'd7268: duty=97; 15'd7269: duty=94; 15'd7270: duty=95; 15'd7271: duty=99;
15'd7272: duty=99; 15'd7273: duty=99; 15'd7274: duty=93; 15'd7275: duty=94; 15'd7276: duty=95; 15'd7277: duty=94; 15'd7278: duty=101; 15'd7279: duty=100;
15'd7280: duty=98; 15'd7281: duty=111; 15'd7282: duty=113; 15'd7283: duty=116; 15'd7284: duty=121; 15'd7285: duty=119; 15'd7286: duty=120; 15'd7287: duty=119;
15'd7288: duty=112; 15'd7289: duty=117; 15'd7290: duty=113; 15'd7291: duty=105; 15'd7292: duty=116; 15'd7293: duty=117; 15'd7294: duty=123; 15'd7295: duty=137;
15'd7296: duty=141; 15'd7297: duty=143; 15'd7298: duty=158; 15'd7299: duty=163; 15'd7300: duty=170; 15'd7301: duty=174; 15'd7302: duty=178; 15'd7303: duty=174;
15'd7304: duty=171; 15'd7305: duty=166; 15'd7306: duty=171; 15'd7307: duty=165; 15'd7308: duty=159; 15'd7309: duty=160; 15'd7310: duty=153; 15'd7311: duty=157;
15'd7312: duty=158; 15'd7313: duty=163; 15'd7314: duty=153; 15'd7315: duty=152; 15'd7316: duty=153; 15'd7317: duty=157; 15'd7318: duty=161; 15'd7319: duty=157;
15'd7320: duty=151; 15'd7321: duty=149; 15'd7322: duty=149; 15'd7323: duty=143; 15'd7324: duty=138; 15'd7325: duty=134; 15'd7326: duty=123; 15'd7327: duty=122;
15'd7328: duty=120; 15'd7329: duty=119; 15'd7330: duty=114; 15'd7331: duty=108; 15'd7332: duty=107; 15'd7333: duty=102; 15'd7334: duty=103; 15'd7335: duty=105;
15'd7336: duty=100; 15'd7337: duty=97; 15'd7338: duty=95; 15'd7339: duty=96; 15'd7340: duty=98; 15'd7341: duty=96; 15'd7342: duty=98; 15'd7343: duty=99;
15'd7344: duty=96; 15'd7345: duty=94; 15'd7346: duty=96; 15'd7347: duty=99; 15'd7348: duty=102; 15'd7349: duty=104; 15'd7350: duty=107; 15'd7351: duty=114;
15'd7352: duty=124; 15'd7353: duty=118; 15'd7354: duty=115; 15'd7355: duty=121; 15'd7356: duty=126; 15'd7357: duty=131; 15'd7358: duty=135; 15'd7359: duty=143;
15'd7360: duty=148; 15'd7361: duty=148; 15'd7362: duty=153; 15'd7363: duty=163; 15'd7364: duty=165; 15'd7365: duty=162; 15'd7366: duty=162; 15'd7367: duty=163;
15'd7368: duty=165; 15'd7369: duty=162; 15'd7370: duty=154; 15'd7371: duty=148; 15'd7372: duty=154; 15'd7373: duty=149; 15'd7374: duty=142; 15'd7375: duty=142;
15'd7376: duty=139; 15'd7377: duty=139; 15'd7378: duty=142; 15'd7379: duty=145; 15'd7380: duty=146; 15'd7381: duty=145; 15'd7382: duty=151; 15'd7383: duty=150;
15'd7384: duty=147; 15'd7385: duty=151; 15'd7386: duty=142; 15'd7387: duty=139; 15'd7388: duty=142; 15'd7389: duty=136; 15'd7390: duty=128; 15'd7391: duty=127;
15'd7392: duty=126; 15'd7393: duty=121; 15'd7394: duty=109; 15'd7395: duty=109; 15'd7396: duty=113; 15'd7397: duty=115; 15'd7398: duty=107; 15'd7399: duty=107;
15'd7400: duty=112; 15'd7401: duty=113; 15'd7402: duty=121; 15'd7403: duty=116; 15'd7404: duty=107; 15'd7405: duty=118; 15'd7406: duty=124; 15'd7407: duty=110;
15'd7408: duty=106; 15'd7409: duty=108; 15'd7410: duty=107; 15'd7411: duty=102; 15'd7412: duty=101; 15'd7413: duty=104; 15'd7414: duty=99; 15'd7415: duty=101;
15'd7416: duty=105; 15'd7417: duty=112; 15'd7418: duty=119; 15'd7419: duty=116; 15'd7420: duty=124; 15'd7421: duty=124; 15'd7422: duty=123; 15'd7423: duty=134;
15'd7424: duty=141; 15'd7425: duty=137; 15'd7426: duty=139; 15'd7427: duty=148; 15'd7428: duty=149; 15'd7429: duty=152; 15'd7430: duty=154; 15'd7431: duty=154;
15'd7432: duty=156; 15'd7433: duty=158; 15'd7434: duty=159; 15'd7435: duty=152; 15'd7436: duty=151; 15'd7437: duty=156; 15'd7438: duty=157; 15'd7439: duty=151;
15'd7440: duty=150; 15'd7441: duty=149; 15'd7442: duty=150; 15'd7443: duty=156; 15'd7444: duty=151; 15'd7445: duty=149; 15'd7446: duty=151; 15'd7447: duty=151;
15'd7448: duty=150; 15'd7449: duty=148; 15'd7450: duty=142; 15'd7451: duty=139; 15'd7452: duty=144; 15'd7453: duty=143; 15'd7454: duty=139; 15'd7455: duty=139;
15'd7456: duty=134; 15'd7457: duty=131; 15'd7458: duty=128; 15'd7459: duty=128; 15'd7460: duty=125; 15'd7461: duty=121; 15'd7462: duty=115; 15'd7463: duty=118;
15'd7464: duty=109; 15'd7465: duty=107; 15'd7466: duty=113; 15'd7467: duty=110; 15'd7468: duty=110; 15'd7469: duty=108; 15'd7470: duty=111; 15'd7471: duty=112;
15'd7472: duty=110; 15'd7473: duty=110; 15'd7474: duty=110; 15'd7475: duty=113; 15'd7476: duty=113; 15'd7477: duty=115; 15'd7478: duty=113; 15'd7479: duty=107;
15'd7480: duty=115; 15'd7481: duty=119; 15'd7482: duty=118; 15'd7483: duty=122; 15'd7484: duty=124; 15'd7485: duty=119; 15'd7486: duty=124; 15'd7487: duty=125;
15'd7488: duty=127; 15'd7489: duty=127; 15'd7490: duty=125; 15'd7491: duty=126; 15'd7492: duty=125; 15'd7493: duty=128; 15'd7494: duty=132; 15'd7495: duty=130;
15'd7496: duty=131; 15'd7497: duty=134; 15'd7498: duty=143; 15'd7499: duty=147; 15'd7500: duty=148; 15'd7501: duty=145; 15'd7502: duty=145; 15'd7503: duty=150;
15'd7504: duty=148; 15'd7505: duty=144; 15'd7506: duty=143; 15'd7507: duty=145; 15'd7508: duty=145; 15'd7509: duty=143; 15'd7510: duty=136; 15'd7511: duty=142;
15'd7512: duty=142; 15'd7513: duty=136; 15'd7514: duty=134; 15'd7515: duty=141; 15'd7516: duty=136; 15'd7517: duty=133; 15'd7518: duty=134; 15'd7519: duty=134;
15'd7520: duty=138; 15'd7521: duty=138; 15'd7522: duty=141; 15'd7523: duty=142; 15'd7524: duty=140; 15'd7525: duty=141; 15'd7526: duty=136; 15'd7527: duty=137;
15'd7528: duty=129; 15'd7529: duty=128; 15'd7530: duty=127; 15'd7531: duty=119; 15'd7532: duty=121; 15'd7533: duty=116; 15'd7534: duty=113; 15'd7535: duty=109;
15'd7536: duty=108; 15'd7537: duty=107; 15'd7538: duty=110; 15'd7539: duty=113; 15'd7540: duty=121; 15'd7541: duty=128; 15'd7542: duty=129; 15'd7543: duty=139;
15'd7544: duty=149; 15'd7545: duty=153; 15'd7546: duty=154; 15'd7547: duty=148; 15'd7548: duty=145; 15'd7549: duty=143; 15'd7550: duty=137; 15'd7551: duty=128;
15'd7552: duty=127; 15'd7553: duty=128; 15'd7554: duty=126; 15'd7555: duty=122; 15'd7556: duty=121; 15'd7557: duty=125; 15'd7558: duty=127; 15'd7559: duty=134;
15'd7560: duty=142; 15'd7561: duty=137; 15'd7562: duty=139; 15'd7563: duty=146; 15'd7564: duty=147; 15'd7565: duty=148; 15'd7566: duty=147; 15'd7567: duty=145;
15'd7568: duty=141; 15'd7569: duty=146; 15'd7570: duty=137; 15'd7571: duty=129; 15'd7572: duty=134; 15'd7573: duty=132; 15'd7574: duty=126; 15'd7575: duty=118;
15'd7576: duty=119; 15'd7577: duty=121; 15'd7578: duty=123; 15'd7579: duty=125; 15'd7580: duty=124; 15'd7581: duty=121; 15'd7582: duty=118; 15'd7583: duty=116;
15'd7584: duty=119; 15'd7585: duty=122; 15'd7586: duty=122; 15'd7587: duty=122; 15'd7588: duty=113; 15'd7589: duty=113; 15'd7590: duty=116; 15'd7591: duty=118;
15'd7592: duty=112; 15'd7593: duty=107; 15'd7594: duty=115; 15'd7595: duty=116; 15'd7596: duty=112; 15'd7597: duty=113; 15'd7598: duty=115; 15'd7599: duty=118;
15'd7600: duty=122; 15'd7601: duty=124; 15'd7602: duty=125; 15'd7603: duty=126; 15'd7604: duty=131; 15'd7605: duty=128; 15'd7606: duty=128; 15'd7607: duty=129;
15'd7608: duty=130; 15'd7609: duty=136; 15'd7610: duty=136; 15'd7611: duty=142; 15'd7612: duty=142; 15'd7613: duty=136; 15'd7614: duty=143; 15'd7615: duty=148;
15'd7616: duty=146; 15'd7617: duty=143; 15'd7618: duty=154; 15'd7619: duty=159; 15'd7620: duty=159; 15'd7621: duty=156; 15'd7622: duty=150; 15'd7623: duty=152;
15'd7624: duty=153; 15'd7625: duty=151; 15'd7626: duty=151; 15'd7627: duty=148; 15'd7628: duty=142; 15'd7629: duty=148; 15'd7630: duty=150; 15'd7631: duty=146;
15'd7632: duty=153; 15'd7633: duty=149; 15'd7634: duty=145; 15'd7635: duty=152; 15'd7636: duty=150; 15'd7637: duty=146; 15'd7638: duty=140; 15'd7639: duty=136;
15'd7640: duty=136; 15'd7641: duty=132; 15'd7642: duty=130; 15'd7643: duty=125; 15'd7644: duty=121; 15'd7645: duty=122; 15'd7646: duty=126; 15'd7647: duty=127;
15'd7648: duty=124; 15'd7649: duty=122; 15'd7650: duty=124; 15'd7651: duty=118; 15'd7652: duty=116; 15'd7653: duty=108; 15'd7654: duty=107; 15'd7655: duty=113;
15'd7656: duty=105; 15'd7657: duty=104; 15'd7658: duty=100; 15'd7659: duty=98; 15'd7660: duty=99; 15'd7661: duty=104; 15'd7662: duty=102; 15'd7663: duty=102;
15'd7664: duty=97; 15'd7665: duty=103; 15'd7666: duty=107; 15'd7667: duty=104; 15'd7668: duty=111; 15'd7669: duty=117; 15'd7670: duty=121; 15'd7671: duty=123;
15'd7672: duty=128; 15'd7673: duty=126; 15'd7674: duty=128; 15'd7675: duty=134; 15'd7676: duty=137; 15'd7677: duty=134; 15'd7678: duty=136; 15'd7679: duty=139;
15'd7680: duty=142; 15'd7681: duty=139; 15'd7682: duty=145; 15'd7683: duty=145; 15'd7684: duty=145; 15'd7685: duty=144; 15'd7686: duty=146; 15'd7687: duty=139;
15'd7688: duty=136; 15'd7689: duty=144; 15'd7690: duty=148; 15'd7691: duty=144; 15'd7692: duty=142; 15'd7693: duty=148; 15'd7694: duty=153; 15'd7695: duty=159;
15'd7696: duty=159; 15'd7697: duty=160; 15'd7698: duty=159; 15'd7699: duty=162; 15'd7700: duty=160; 15'd7701: duty=160; 15'd7702: duty=153; 15'd7703: duty=148;
15'd7704: duty=142; 15'd7705: duty=142; 15'd7706: duty=139; 15'd7707: duty=134; 15'd7708: duty=133; 15'd7709: duty=130; 15'd7710: duty=125; 15'd7711: duty=128;
15'd7712: duty=129; 15'd7713: duty=124; 15'd7714: duty=125; 15'd7715: duty=125; 15'd7716: duty=127; 15'd7717: duty=125; 15'd7718: duty=121; 15'd7719: duty=124;
15'd7720: duty=127; 15'd7721: duty=124; 15'd7722: duty=119; 15'd7723: duty=112; 15'd7724: duty=109; 15'd7725: duty=107; 15'd7726: duty=107; 15'd7727: duty=107;
15'd7728: duty=108; 15'd7729: duty=107; 15'd7730: duty=105; 15'd7731: duty=105; 15'd7732: duty=108; 15'd7733: duty=109; 15'd7734: duty=114; 15'd7735: duty=113;
15'd7736: duty=119; 15'd7737: duty=122; 15'd7738: duty=119; 15'd7739: duty=123; 15'd7740: duty=124; 15'd7741: duty=130; 15'd7742: duty=131; 15'd7743: duty=136;
15'd7744: duty=134; 15'd7745: duty=134; 15'd7746: duty=137; 15'd7747: duty=139; 15'd7748: duty=136; 15'd7749: duty=137; 15'd7750: duty=142; 15'd7751: duty=143;
15'd7752: duty=137; 15'd7753: duty=137; 15'd7754: duty=143; 15'd7755: duty=140; 15'd7756: duty=140; 15'd7757: duty=147; 15'd7758: duty=145; 15'd7759: duty=145;
15'd7760: duty=151; 15'd7761: duty=150; 15'd7762: duty=153; 15'd7763: duty=154; 15'd7764: duty=156; 15'd7765: duty=156; 15'd7766: duty=152; 15'd7767: duty=145;
15'd7768: duty=149; 15'd7769: duty=144; 15'd7770: duty=139; 15'd7771: duty=140; 15'd7772: duty=139; 15'd7773: duty=134; 15'd7774: duty=130; 15'd7775: duty=136;
15'd7776: duty=136; 15'd7777: duty=131; 15'd7778: duty=125; 15'd7779: duty=125; 15'd7780: duty=128; 15'd7781: duty=129; 15'd7782: duty=122; 15'd7783: duty=124;
15'd7784: duty=122; 15'd7785: duty=119; 15'd7786: duty=125; 15'd7787: duty=122; 15'd7788: duty=113; 15'd7789: duty=112; 15'd7790: duty=116; 15'd7791: duty=111;
15'd7792: duty=107; 15'd7793: duty=110; 15'd7794: duty=113; 15'd7795: duty=113; 15'd7796: duty=107; 15'd7797: duty=107; 15'd7798: duty=107; 15'd7799: duty=105;
15'd7800: duty=99; 15'd7801: duty=104; 15'd7802: duty=110; 15'd7803: duty=111; 15'd7804: duty=123; 15'd7805: duty=128; 15'd7806: duty=131; 15'd7807: duty=134;
15'd7808: duty=138; 15'd7809: duty=140; 15'd7810: duty=142; 15'd7811: duty=142; 15'd7812: duty=138; 15'd7813: duty=135; 15'd7814: duty=133; 15'd7815: duty=135;
15'd7816: duty=134; 15'd7817: duty=138; 15'd7818: duty=137; 15'd7819: duty=137; 15'd7820: duty=148; 15'd7821: duty=154; 15'd7822: duty=154; 15'd7823: duty=154;
15'd7824: duty=154; 15'd7825: duty=155; 15'd7826: duty=157; 15'd7827: duty=149; 15'd7828: duty=148; 15'd7829: duty=148; 15'd7830: duty=144; 15'd7831: duty=142;
15'd7832: duty=140; 15'd7833: duty=138; 15'd7834: duty=137; 15'd7835: duty=136; 15'd7836: duty=134; 15'd7837: duty=137; 15'd7838: duty=134; 15'd7839: duty=134;
15'd7840: duty=133; 15'd7841: duty=136; 15'd7842: duty=133; 15'd7843: duty=129; 15'd7844: duty=133; 15'd7845: duty=129; 15'd7846: duty=126; 15'd7847: duty=118;
15'd7848: duty=115; 15'd7849: duty=119; 15'd7850: duty=118; 15'd7851: duty=117; 15'd7852: duty=119; 15'd7853: duty=119; 15'd7854: duty=121; 15'd7855: duty=119;
15'd7856: duty=117; 15'd7857: duty=122; 15'd7858: duty=124; 15'd7859: duty=119; 15'd7860: duty=120; 15'd7861: duty=128; 15'd7862: duty=124; 15'd7863: duty=124;
15'd7864: duty=123; 15'd7865: duty=125; 15'd7866: duty=128; 15'd7867: duty=127; 15'd7868: duty=127; 15'd7869: duty=131; 15'd7870: duty=133; 15'd7871: duty=133;
15'd7872: duty=136; 15'd7873: duty=134; 15'd7874: duty=134; 15'd7875: duty=134; 15'd7876: duty=136; 15'd7877: duty=134; 15'd7878: duty=133; 15'd7879: duty=128;
15'd7880: duty=126; 15'd7881: duty=122; 15'd7882: duty=124; 15'd7883: duty=124; 15'd7884: duty=120; 15'd7885: duty=125; 15'd7886: duty=128; 15'd7887: duty=129;
15'd7888: duty=130; 15'd7889: duty=139; 15'd7890: duty=137; 15'd7891: duty=135; 15'd7892: duty=136; 15'd7893: duty=140; 15'd7894: duty=141; 15'd7895: duty=138;
15'd7896: duty=137; 15'd7897: duty=140; 15'd7898: duty=137; 15'd7899: duty=134; 15'd7900: duty=134; 15'd7901: duty=132; 15'd7902: duty=127; 15'd7903: duty=124;
15'd7904: duty=130; 15'd7905: duty=125; 15'd7906: duty=125; 15'd7907: duty=128; 15'd7908: duty=131; 15'd7909: duty=134; 15'd7910: duty=131; 15'd7911: duty=134;
15'd7912: duty=133; 15'd7913: duty=130; 15'd7914: duty=126; 15'd7915: duty=125; 15'd7916: duty=120; 15'd7917: duty=115; 15'd7918: duty=112; 15'd7919: duty=105;
15'd7920: duty=109; 15'd7921: duty=111; 15'd7922: duty=113; 15'd7923: duty=119; 15'd7924: duty=123; 15'd7925: duty=128; 15'd7926: duty=128; 15'd7927: duty=127;
15'd7928: duty=128; 15'd7929: duty=130; 15'd7930: duty=136; 15'd7931: duty=136; 15'd7932: duty=131; 15'd7933: duty=133; 15'd7934: duty=138; 15'd7935: duty=134;
15'd7936: duty=130; 15'd7937: duty=133; 15'd7938: duty=139; 15'd7939: duty=143; 15'd7940: duty=142; 15'd7941: duty=140; 15'd7942: duty=141; 15'd7943: duty=140;
15'd7944: duty=147; 15'd7945: duty=149; 15'd7946: duty=145; 15'd7947: duty=143; 15'd7948: duty=147; 15'd7949: duty=148; 15'd7950: duty=142; 15'd7951: duty=138;
15'd7952: duty=139; 15'd7953: duty=140; 15'd7954: duty=138; 15'd7955: duty=137; 15'd7956: duty=137; 15'd7957: duty=140; 15'd7958: duty=147; 15'd7959: duty=152;
15'd7960: duty=151; 15'd7961: duty=148; 15'd7962: duty=147; 15'd7963: duty=143; 15'd7964: duty=139; 15'd7965: duty=139; 15'd7966: duty=133; 15'd7967: duty=131;
15'd7968: duty=127; 15'd7969: duty=132; 15'd7970: duty=126; 15'd7971: duty=119; 15'd7972: duty=124; 15'd7973: duty=128; 15'd7974: duty=124; 15'd7975: duty=122;
15'd7976: duty=124; 15'd7977: duty=128; 15'd7978: duty=121; 15'd7979: duty=122; 15'd7980: duty=124; 15'd7981: duty=117; 15'd7982: duty=115; 15'd7983: duty=113;
15'd7984: duty=112; 15'd7985: duty=109; 15'd7986: duty=107; 15'd7987: duty=105; 15'd7988: duty=109; 15'd7989: duty=107; 15'd7990: duty=112; 15'd7991: duty=115;
15'd7992: duty=110; 15'd7993: duty=110; 15'd7994: duty=117; 15'd7995: duty=116; 15'd7996: duty=115; 15'd7997: duty=118; 15'd7998: duty=118; 15'd7999: duty=119;
15'd8000: duty=121; 15'd8001: duty=122; 15'd8002: duty=123; 15'd8003: duty=118; 15'd8004: duty=121; 15'd8005: duty=127; 15'd8006: duty=127; 15'd8007: duty=124;
15'd8008: duty=128; 15'd8009: duty=132; 15'd8010: duty=130; 15'd8011: duty=132; 15'd8012: duty=134; 15'd8013: duty=135; 15'd8014: duty=134; 15'd8015: duty=137;
15'd8016: duty=138; 15'd8017: duty=137; 15'd8018: duty=139; 15'd8019: duty=140; 15'd8020: duty=142; 15'd8021: duty=146; 15'd8022: duty=144; 15'd8023: duty=148;
15'd8024: duty=153; 15'd8025: duty=153; 15'd8026: duty=154; 15'd8027: duty=156; 15'd8028: duty=153; 15'd8029: duty=150; 15'd8030: duty=150; 15'd8031: duty=151;
15'd8032: duty=150; 15'd8033: duty=140; 15'd8034: duty=136; 15'd8035: duty=140; 15'd8036: duty=142; 15'd8037: duty=137; 15'd8038: duty=141; 15'd8039: duty=140;
15'd8040: duty=139; 15'd8041: duty=145; 15'd8042: duty=144; 15'd8043: duty=140; 15'd8044: duty=131; 15'd8045: duty=134; 15'd8046: duty=134; 15'd8047: duty=128;
15'd8048: duty=127; 15'd8049: duty=125; 15'd8050: duty=124; 15'd8051: duty=127; 15'd8052: duty=127; 15'd8053: duty=125; 15'd8054: duty=126; 15'd8055: duty=127;
15'd8056: duty=122; 15'd8057: duty=119; 15'd8058: duty=125; 15'd8059: duty=127; 15'd8060: duty=121; 15'd8061: duty=124; 15'd8062: duty=128; 15'd8063: duty=124;
15'd8064: duty=124; 15'd8065: duty=125; 15'd8066: duty=126; 15'd8067: duty=124; 15'd8068: duty=122; 15'd8069: duty=118; 15'd8070: duty=118; 15'd8071: duty=118;
15'd8072: duty=119; 15'd8073: duty=121; 15'd8074: duty=119; 15'd8075: duty=118; 15'd8076: duty=124; 15'd8077: duty=130; 15'd8078: duty=131; 15'd8079: duty=128;
15'd8080: duty=127; 15'd8081: duty=128; 15'd8082: duty=134; 15'd8083: duty=131; 15'd8084: duty=127; 15'd8085: duty=131; 15'd8086: duty=131; 15'd8087: duty=134;
15'd8088: duty=137; 15'd8089: duty=137; 15'd8090: duty=137; 15'd8091: duty=140; 15'd8092: duty=136; 15'd8093: duty=139; 15'd8094: duty=140; 15'd8095: duty=136;
15'd8096: duty=134; 15'd8097: duty=139; 15'd8098: duty=136; 15'd8099: duty=130; 15'd8100: duty=131; 15'd8101: duty=131; 15'd8102: duty=131; 15'd8103: duty=127;
15'd8104: duty=124; 15'd8105: duty=127; 15'd8106: duty=128; 15'd8107: duty=124; 15'd8108: duty=124; 15'd8109: duty=131; 15'd8110: duty=133; 15'd8111: duty=130;
15'd8112: duty=127; 15'd8113: duty=128; 15'd8114: duty=132; 15'd8115: duty=130; 15'd8116: duty=127; 15'd8117: duty=130; 15'd8118: duty=131; 15'd8119: duty=128;
15'd8120: duty=128; 15'd8121: duty=124; 15'd8122: duty=122; 15'd8123: duty=125; 15'd8124: duty=124; 15'd8125: duty=122; 15'd8126: duty=124; 15'd8127: duty=124;
15'd8128: duty=124; 15'd8129: duty=127; 15'd8130: duty=127; 15'd8131: duty=126; 15'd8132: duty=130; 15'd8133: duty=133; 15'd8134: duty=137; 15'd8135: duty=139;
15'd8136: duty=137; 15'd8137: duty=133; 15'd8138: duty=133; 15'd8139: duty=133; 15'd8140: duty=134; 15'd8141: duty=131; 15'd8142: duty=133; 15'd8143: duty=134;
15'd8144: duty=134; 15'd8145: duty=136; 15'd8146: duty=139; 15'd8147: duty=134; 15'd8148: duty=129; 15'd8149: duty=134; 15'd8150: duty=139; 15'd8151: duty=140;
15'd8152: duty=137; 15'd8153: duty=133; 15'd8154: duty=136; 15'd8155: duty=137; 15'd8156: duty=136; 15'd8157: duty=139; 15'd8158: duty=136; 15'd8159: duty=134;
15'd8160: duty=136; 15'd8161: duty=139; 15'd8162: duty=136; 15'd8163: duty=134; 15'd8164: duty=133; 15'd8165: duty=133; 15'd8166: duty=127; 15'd8167: duty=128;
15'd8168: duty=127; 15'd8169: duty=128; 15'd8170: duty=128; 15'd8171: duty=126; 15'd8172: duty=128; 15'd8173: duty=124; 15'd8174: duty=119; 15'd8175: duty=122;
15'd8176: duty=125; 15'd8177: duty=127; 15'd8178: duty=129; 15'd8179: duty=130; 15'd8180: duty=134; 15'd8181: duty=133; 15'd8182: duty=131; 15'd8183: duty=137;
15'd8184: duty=139; 15'd8185: duty=131; 15'd8186: duty=137; 15'd8187: duty=139; 15'd8188: duty=134; 15'd8189: duty=133; 15'd8190: duty=137; 15'd8191: duty=133;
15'd8192: duty=132; 15'd8193: duty=133; 15'd8194: duty=131; 15'd8195: duty=133; 15'd8196: duty=134; 15'd8197: duty=131; 15'd8198: duty=131; 15'd8199: duty=133;
15'd8200: duty=128; 15'd8201: duty=127; 15'd8202: duty=132; 15'd8203: duty=130; 15'd8204: duty=125; 15'd8205: duty=124; 15'd8206: duty=124; 15'd8207: duty=124;
15'd8208: duty=127; 15'd8209: duty=126; 15'd8210: duty=127; 15'd8211: duty=131; 15'd8212: duty=136; 15'd8213: duty=134; 15'd8214: duty=132; 15'd8215: duty=131;
15'd8216: duty=131; 15'd8217: duty=134; 15'd8218: duty=136; 15'd8219: duty=133; 15'd8220: duty=121; 15'd8221: duty=118; 15'd8222: duty=121; 15'd8223: duty=121;
15'd8224: duty=119; 15'd8225: duty=119; 15'd8226: duty=116; 15'd8227: duty=119; 15'd8228: duty=126; 15'd8229: duty=127; 15'd8230: duty=127; 15'd8231: duty=125;
15'd8232: duty=124; 15'd8233: duty=129; 15'd8234: duty=128; 15'd8235: duty=124; 15'd8236: duty=121; 15'd8237: duty=127; 15'd8238: duty=126; 15'd8239: duty=122;
15'd8240: duty=121; 15'd8241: duty=117; 15'd8242: duty=116; 15'd8243: duty=124; 15'd8244: duty=124; 15'd8245: duty=119; 15'd8246: duty=121; 15'd8247: duty=125;
15'd8248: duty=124; 15'd8249: duty=128; 15'd8250: duty=127; 15'd8251: duty=134; 15'd8252: duty=137; 15'd8253: duty=134; 15'd8254: duty=141; 15'd8255: duty=143;
15'd8256: duty=147; 15'd8257: duty=145; 15'd8258: duty=145; 15'd8259: duty=145; 15'd8260: duty=144; 15'd8261: duty=142; 15'd8262: duty=144; 15'd8263: duty=143;
15'd8264: duty=142; 15'd8265: duty=146; 15'd8266: duty=147; 15'd8267: duty=149; 15'd8268: duty=148; 15'd8269: duty=148; 15'd8270: duty=147; 15'd8271: duty=148;
15'd8272: duty=147; 15'd8273: duty=145; 15'd8274: duty=147; 15'd8275: duty=149; 15'd8276: duty=151; 15'd8277: duty=145; 15'd8278: duty=138; 15'd8279: duty=145;
15'd8280: duty=144; 15'd8281: duty=140; 15'd8282: duty=137; 15'd8283: duty=135; 15'd8284: duty=131; 15'd8285: duty=131; 15'd8286: duty=130; 15'd8287: duty=125;
15'd8288: duty=123; 15'd8289: duty=119; 15'd8290: duty=118; 15'd8291: duty=124; 15'd8292: duty=120; 15'd8293: duty=118; 15'd8294: duty=117; 15'd8295: duty=116;
15'd8296: duty=118; 15'd8297: duty=122; 15'd8298: duty=120; 15'd8299: duty=119; 15'd8300: duty=121; 15'd8301: duty=119; 15'd8302: duty=118; 15'd8303: duty=112;
15'd8304: duty=110; 15'd8305: duty=107; 15'd8306: duty=113; 15'd8307: duty=111; 15'd8308: duty=110; 15'd8309: duty=110; 15'd8310: duty=110; 15'd8311: duty=118;
15'd8312: duty=119; 15'd8313: duty=119; 15'd8314: duty=124; 15'd8315: duty=119; 15'd8316: duty=121; 15'd8317: duty=128; 15'd8318: duty=125; 15'd8319: duty=124;
15'd8320: duty=128; 15'd8321: duty=133; 15'd8322: duty=133; 15'd8323: duty=137; 15'd8324: duty=136; 15'd8325: duty=133; 15'd8326: duty=131; 15'd8327: duty=134;
15'd8328: duty=134; 15'd8329: duty=134; 15'd8330: duty=134; 15'd8331: duty=139; 15'd8332: duty=142; 15'd8333: duty=141; 15'd8334: duty=139; 15'd8335: duty=140;
15'd8336: duty=148; 15'd8337: duty=148; 15'd8338: duty=143; 15'd8339: duty=143; 15'd8340: duty=146; 15'd8341: duty=141; 15'd8342: duty=143; 15'd8343: duty=144;
15'd8344: duty=139; 15'd8345: duty=137; 15'd8346: duty=136; 15'd8347: duty=137; 15'd8348: duty=143; 15'd8349: duty=137; 15'd8350: duty=131; 15'd8351: duty=133;
15'd8352: duty=133; 15'd8353: duty=129; 15'd8354: duty=127; 15'd8355: duty=131; 15'd8356: duty=127; 15'd8357: duty=127; 15'd8358: duty=126; 15'd8359: duty=124;
15'd8360: duty=122; 15'd8361: duty=118; 15'd8362: duty=115; 15'd8363: duty=118; 15'd8364: duty=122; 15'd8365: duty=119; 15'd8366: duty=123; 15'd8367: duty=119;
15'd8368: duty=121; 15'd8369: duty=128; 15'd8370: duty=128; 15'd8371: duty=135; 15'd8372: duty=133; 15'd8373: duty=134; 15'd8374: duty=136; 15'd8375: duty=129;
15'd8376: duty=124; 15'd8377: duty=132; 15'd8378: duty=134; 15'd8379: duty=137; 15'd8380: duty=142; 15'd8381: duty=140; 15'd8382: duty=142; 15'd8383: duty=142;
15'd8384: duty=138; 15'd8385: duty=136; 15'd8386: duty=142; 15'd8387: duty=142; 15'd8388: duty=141; 15'd8389: duty=143; 15'd8390: duty=145; 15'd8391: duty=145;
15'd8392: duty=142; 15'd8393: duty=140; 15'd8394: duty=144; 15'd8395: duty=143; 15'd8396: duty=139; 15'd8397: duty=139; 15'd8398: duty=140; 15'd8399: duty=140;
15'd8400: duty=136; 15'd8401: duty=134; 15'd8402: duty=136; 15'd8403: duty=133; 15'd8404: duty=128; 15'd8405: duty=130; 15'd8406: duty=131; 15'd8407: duty=127;
15'd8408: duty=124; 15'd8409: duty=124; 15'd8410: duty=119; 15'd8411: duty=115; 15'd8412: duty=118; 15'd8413: duty=115; 15'd8414: duty=113; 15'd8415: duty=113;
15'd8416: duty=113; 15'd8417: duty=112; 15'd8418: duty=112; 15'd8419: duty=110; 15'd8420: duty=115; 15'd8421: duty=115; 15'd8422: duty=112; 15'd8423: duty=112;
15'd8424: duty=107; 15'd8425: duty=112; 15'd8426: duty=112; 15'd8427: duty=110; 15'd8428: duty=110; 15'd8429: duty=107; 15'd8430: duty=105; 15'd8431: duty=104;
15'd8432: duty=102; 15'd8433: duty=105; 15'd8434: duty=108; 15'd8435: duty=110; 15'd8436: duty=118; 15'd8437: duty=124; 15'd8438: duty=129; 15'd8439: duty=134;
15'd8440: duty=139; 15'd8441: duty=142; 15'd8442: duty=153; 15'd8443: duty=153; 15'd8444: duty=145; 15'd8445: duty=143; 15'd8446: duty=146; 15'd8447: duty=146;
15'd8448: duty=145; 15'd8449: duty=143; 15'd8450: duty=136; 15'd8451: duty=144; 15'd8452: duty=150; 15'd8453: duty=156; 15'd8454: duty=156; 15'd8455: duty=154;
15'd8456: duty=159; 15'd8457: duty=163; 15'd8458: duty=162; 15'd8459: duty=160; 15'd8460: duty=160; 15'd8461: duty=160; 15'd8462: duty=162; 15'd8463: duty=159;
15'd8464: duty=153; 15'd8465: duty=146; 15'd8466: duty=145; 15'd8467: duty=146; 15'd8468: duty=148; 15'd8469: duty=146; 15'd8470: duty=143; 15'd8471: duty=148;
15'd8472: duty=148; 15'd8473: duty=148; 15'd8474: duty=144; 15'd8475: duty=139; 15'd8476: duty=139; 15'd8477: duty=142; 15'd8478: duty=136; 15'd8479: duty=128;
15'd8480: duty=126; 15'd8481: duty=118; 15'd8482: duty=116; 15'd8483: duty=118; 15'd8484: duty=115; 15'd8485: duty=111; 15'd8486: duty=106; 15'd8487: duty=108;
15'd8488: duty=115; 15'd8489: duty=113; 15'd8490: duty=107; 15'd8491: duty=107; 15'd8492: duty=112; 15'd8493: duty=108; 15'd8494: duty=106; 15'd8495: duty=104;
15'd8496: duty=104; 15'd8497: duty=104; 15'd8498: duty=104; 15'd8499: duty=104; 15'd8500: duty=104; 15'd8501: duty=102; 15'd8502: duty=101; 15'd8503: duty=108;
15'd8504: duty=107; 15'd8505: duty=108; 15'd8506: duty=112; 15'd8507: duty=113; 15'd8508: duty=112; 15'd8509: duty=118; 15'd8510: duty=124; 15'd8511: duty=126;
15'd8512: duty=125; 15'd8513: duty=128; 15'd8514: duty=134; 15'd8515: duty=139; 15'd8516: duty=137; 15'd8517: duty=137; 15'd8518: duty=139; 15'd8519: duty=142;
15'd8520: duty=146; 15'd8521: duty=148; 15'd8522: duty=143; 15'd8523: duty=145; 15'd8524: duty=149; 15'd8525: duty=148; 15'd8526: duty=149; 15'd8527: duty=150;
15'd8528: duty=151; 15'd8529: duty=157; 15'd8530: duty=160; 15'd8531: duty=158; 15'd8532: duty=156; 15'd8533: duty=153; 15'd8534: duty=151; 15'd8535: duty=154;
15'd8536: duty=153; 15'd8537: duty=147; 15'd8538: duty=142; 15'd8539: duty=144; 15'd8540: duty=146; 15'd8541: duty=143; 15'd8542: duty=145; 15'd8543: duty=139;
15'd8544: duty=137; 15'd8545: duty=136; 15'd8546: duty=133; 15'd8547: duty=130; 15'd8548: duty=127; 15'd8549: duty=127; 15'd8550: duty=130; 15'd8551: duty=127;
15'd8552: duty=122; 15'd8553: duty=119; 15'd8554: duty=118; 15'd8555: duty=118; 15'd8556: duty=119; 15'd8557: duty=119; 15'd8558: duty=115; 15'd8559: duty=114;
15'd8560: duty=116; 15'd8561: duty=118; 15'd8562: duty=118; 15'd8563: duty=116; 15'd8564: duty=110; 15'd8565: duty=113; 15'd8566: duty=116; 15'd8567: duty=116;
15'd8568: duty=118; 15'd8569: duty=116; 15'd8570: duty=115; 15'd8571: duty=119; 15'd8572: duty=126; 15'd8573: duty=122; 15'd8574: duty=127; 15'd8575: duty=132;
15'd8576: duty=130; 15'd8577: duty=137; 15'd8578: duty=138; 15'd8579: duty=131; 15'd8580: duty=133; 15'd8581: duty=136; 15'd8582: duty=131; 15'd8583: duty=132;
15'd8584: duty=130; 15'd8585: duty=131; 15'd8586: duty=134; 15'd8587: duty=135; 15'd8588: duty=133; 15'd8589: duty=134; 15'd8590: duty=134; 15'd8591: duty=135;
15'd8592: duty=136; 15'd8593: duty=139; 15'd8594: duty=142; 15'd8595: duty=142; 15'd8596: duty=141; 15'd8597: duty=139; 15'd8598: duty=142; 15'd8599: duty=140;
15'd8600: duty=142; 15'd8601: duty=140; 15'd8602: duty=140; 15'd8603: duty=140; 15'd8604: duty=142; 15'd8605: duty=137; 15'd8606: duty=137; 15'd8607: duty=139;
15'd8608: duty=139; 15'd8609: duty=137; 15'd8610: duty=131; 15'd8611: duty=128; 15'd8612: duty=126; 15'd8613: duty=124; 15'd8614: duty=122; 15'd8615: duty=122;
15'd8616: duty=122; 15'd8617: duty=116; 15'd8618: duty=118; 15'd8619: duty=121; 15'd8620: duty=118; 15'd8621: duty=116; 15'd8622: duty=115; 15'd8623: duty=113;
15'd8624: duty=118; 15'd8625: duty=124; 15'd8626: duty=118; 15'd8627: duty=116; 15'd8628: duty=118; 15'd8629: duty=125; 15'd8630: duty=125; 15'd8631: duty=119;
15'd8632: duty=119; 15'd8633: duty=118; 15'd8634: duty=121; 15'd8635: duty=127; 15'd8636: duty=127; 15'd8637: duty=125; 15'd8638: duty=125; 15'd8639: duty=130;
15'd8640: duty=133; 15'd8641: duty=136; 15'd8642: duty=133; 15'd8643: duty=130; 15'd8644: duty=136; 15'd8645: duty=142; 15'd8646: duty=142; 15'd8647: duty=143;
15'd8648: duty=142; 15'd8649: duty=145; 15'd8650: duty=151; 15'd8651: duty=154; 15'd8652: duty=148; 15'd8653: duty=148; 15'd8654: duty=150; 15'd8655: duty=150;
15'd8656: duty=154; 15'd8657: duty=148; 15'd8658: duty=142; 15'd8659: duty=143; 15'd8660: duty=145; 15'd8661: duty=145; 15'd8662: duty=144; 15'd8663: duty=142;
15'd8664: duty=140; 15'd8665: duty=137; 15'd8666: duty=142; 15'd8667: duty=137; 15'd8668: duty=128; 15'd8669: duty=131; 15'd8670: duty=133; 15'd8671: duty=131;
15'd8672: duty=131; 15'd8673: duty=128; 15'd8674: duty=126; 15'd8675: duty=125; 15'd8676: duty=126; 15'd8677: duty=127; 15'd8678: duty=125; 15'd8679: duty=121;
15'd8680: duty=119; 15'd8681: duty=121; 15'd8682: duty=121; 15'd8683: duty=122; 15'd8684: duty=116; 15'd8685: duty=112; 15'd8686: duty=115; 15'd8687: duty=115;
15'd8688: duty=118; 15'd8689: duty=118; 15'd8690: duty=113; 15'd8691: duty=112; 15'd8692: duty=117; 15'd8693: duty=119; 15'd8694: duty=118; 15'd8695: duty=115;
15'd8696: duty=119; 15'd8697: duty=121; 15'd8698: duty=122; 15'd8699: duty=124; 15'd8700: duty=121; 15'd8701: duty=118; 15'd8702: duty=122; 15'd8703: duty=127;
15'd8704: duty=125; 15'd8705: duty=126; 15'd8706: duty=127; 15'd8707: duty=131; 15'd8708: duty=131; 15'd8709: duty=135; 15'd8710: duty=131; 15'd8711: duty=131;
15'd8712: duty=130; 15'd8713: duty=136; 15'd8714: duty=145; 15'd8715: duty=141; 15'd8716: duty=137; 15'd8717: duty=137; 15'd8718: duty=140; 15'd8719: duty=141;
15'd8720: duty=146; 15'd8721: duty=141; 15'd8722: duty=142; 15'd8723: duty=144; 15'd8724: duty=140; 15'd8725: duty=137; 15'd8726: duty=134; 15'd8727: duty=133;
15'd8728: duty=138; 15'd8729: duty=142; 15'd8730: duty=142; 15'd8731: duty=142; 15'd8732: duty=146; 15'd8733: duty=144; 15'd8734: duty=143; 15'd8735: duty=145;
15'd8736: duty=142; 15'd8737: duty=134; 15'd8738: duty=131; 15'd8739: duty=134; 15'd8740: duty=134; 15'd8741: duty=128; 15'd8742: duty=127; 15'd8743: duty=128;
15'd8744: duty=128; 15'd8745: duty=134; 15'd8746: duty=131; 15'd8747: duty=127; 15'd8748: duty=130; 15'd8749: duty=128; 15'd8750: duty=129; 15'd8751: duty=126;
15'd8752: duty=125; 15'd8753: duty=126; 15'd8754: duty=120; 15'd8755: duty=124; 15'd8756: duty=131; 15'd8757: duty=121; 15'd8758: duty=119; 15'd8759: duty=124;
15'd8760: duty=122; 15'd8761: duty=123; 15'd8762: duty=121; 15'd8763: duty=121; 15'd8764: duty=121; 15'd8765: duty=121; 15'd8766: duty=134; 15'd8767: duty=131;
15'd8768: duty=125; 15'd8769: duty=125; 15'd8770: duty=127; 15'd8771: duty=130; 15'd8772: duty=131; 15'd8773: duty=128; 15'd8774: duty=127; 15'd8775: duty=128;
15'd8776: duty=131; 15'd8777: duty=136; 15'd8778: duty=132; 15'd8779: duty=131; 15'd8780: duty=129; 15'd8781: duty=131; 15'd8782: duty=137; 15'd8783: duty=137;
15'd8784: duty=136; 15'd8785: duty=140; 15'd8786: duty=140; 15'd8787: duty=140; 15'd8788: duty=136; 15'd8789: duty=133; 15'd8790: duty=138; 15'd8791: duty=133;
15'd8792: duty=134; 15'd8793: duty=137; 15'd8794: duty=128; 15'd8795: duty=124; 15'd8796: duty=127; 15'd8797: duty=130; 15'd8798: duty=128; 15'd8799: duty=123;
15'd8800: duty=129; 15'd8801: duty=131; 15'd8802: duty=129; 15'd8803: duty=134; 15'd8804: duty=134; 15'd8805: duty=128; 15'd8806: duty=132; 15'd8807: duty=130;
15'd8808: duty=131; 15'd8809: duty=133; 15'd8810: duty=129; 15'd8811: duty=130; 15'd8812: duty=128; 15'd8813: duty=131; 15'd8814: duty=128; 15'd8815: duty=123;
15'd8816: duty=124; 15'd8817: duty=121; 15'd8818: duty=127; 15'd8819: duty=136; 15'd8820: duty=139; 15'd8821: duty=131; 15'd8822: duty=132; 15'd8823: duty=139;
15'd8824: duty=134; 15'd8825: duty=137; 15'd8826: duty=136; 15'd8827: duty=133; 15'd8828: duty=136; 15'd8829: duty=143; 15'd8830: duty=140; 15'd8831: duty=134;
15'd8832: duty=131; 15'd8833: duty=128; 15'd8834: duty=134; 15'd8835: duty=139; 15'd8836: duty=134; 15'd8837: duty=128; 15'd8838: duty=127; 15'd8839: duty=135;
15'd8840: duty=136; 15'd8841: duty=133; 15'd8842: duty=131; 15'd8843: duty=129; 15'd8844: duty=136; 15'd8845: duty=137; 15'd8846: duty=130; 15'd8847: duty=125;
15'd8848: duty=120; 15'd8849: duty=121; 15'd8850: duty=124; 15'd8851: duty=125; 15'd8852: duty=122; 15'd8853: duty=117; 15'd8854: duty=122; 15'd8855: duty=123;
15'd8856: duty=123; 15'd8857: duty=118; 15'd8858: duty=121; 15'd8859: duty=125; 15'd8860: duty=128; 15'd8861: duty=134; 15'd8862: duty=130; 15'd8863: duty=128;
15'd8864: duty=133; 15'd8865: duty=131; 15'd8866: duty=130; 15'd8867: duty=129; 15'd8868: duty=127; 15'd8869: duty=129; 15'd8870: duty=128; 15'd8871: duty=127;
15'd8872: duty=128; 15'd8873: duty=131; 15'd8874: duty=130; 15'd8875: duty=131; 15'd8876: duty=135; 15'd8877: duty=131; 15'd8878: duty=130; 15'd8879: duty=132;
15'd8880: duty=131; 15'd8881: duty=128; 15'd8882: duty=134; 15'd8883: duty=131; 15'd8884: duty=128; 15'd8885: duty=136; 15'd8886: duty=136; 15'd8887: duty=137;
15'd8888: duty=130; 15'd8889: duty=137; 15'd8890: duty=139; 15'd8891: duty=129; 15'd8892: duty=134; 15'd8893: duty=140; 15'd8894: duty=136; 15'd8895: duty=131;
15'd8896: duty=133; 15'd8897: duty=137; 15'd8898: duty=139; 15'd8899: duty=137; 15'd8900: duty=130; 15'd8901: duty=134; 15'd8902: duty=136; 15'd8903: duty=136;
15'd8904: duty=138; 15'd8905: duty=129; 15'd8906: duty=130; 15'd8907: duty=128; 15'd8908: duty=131; 15'd8909: duty=129; 15'd8910: duty=126; 15'd8911: duty=131;
15'd8912: duty=130; 15'd8913: duty=129; 15'd8914: duty=128; 15'd8915: duty=129; 15'd8916: duty=128; 15'd8917: duty=131; 15'd8918: duty=131; 15'd8919: duty=129;
15'd8920: duty=133; 15'd8921: duty=128; 15'd8922: duty=123; 15'd8923: duty=125; 15'd8924: duty=128; 15'd8925: duty=122; 15'd8926: duty=115; 15'd8927: duty=114;
15'd8928: duty=110; 15'd8929: duty=117; 15'd8930: duty=120; 15'd8931: duty=122; 15'd8932: duty=121; 15'd8933: duty=127; 15'd8934: duty=135; 15'd8935: duty=141;
15'd8936: duty=135; 15'd8937: duty=132; 15'd8938: duty=139; 15'd8939: duty=131; 15'd8940: duty=130; 15'd8941: duty=129; 15'd8942: duty=130; 15'd8943: duty=128;
15'd8944: duty=130; 15'd8945: duty=129; 15'd8946: duty=131; 15'd8947: duty=137; 15'd8948: duty=137; 15'd8949: duty=137; 15'd8950: duty=134; 15'd8951: duty=143;
15'd8952: duty=142; 15'd8953: duty=145; 15'd8954: duty=145; 15'd8955: duty=139; 15'd8956: duty=136; 15'd8957: duty=133; 15'd8958: duty=139; 15'd8959: duty=137;
15'd8960: duty=136; 15'd8961: duty=134; 15'd8962: duty=133; 15'd8963: duty=136; 15'd8964: duty=131; 15'd8965: duty=132; 15'd8966: duty=139; 15'd8967: duty=134;
15'd8968: duty=130; 15'd8969: duty=127; 15'd8970: duty=128; 15'd8971: duty=129; 15'd8972: duty=128; 15'd8973: duty=134; 15'd8974: duty=136; 15'd8975: duty=140;
15'd8976: duty=137; 15'd8977: duty=133; 15'd8978: duty=133; 15'd8979: duty=127; 15'd8980: duty=126; 15'd8981: duty=122; 15'd8982: duty=121; 15'd8983: duty=126;
15'd8984: duty=118; 15'd8985: duty=116; 15'd8986: duty=127; 15'd8987: duty=128; 15'd8988: duty=128; 15'd8989: duty=124; 15'd8990: duty=116; 15'd8991: duty=119;
15'd8992: duty=127; 15'd8993: duty=124; 15'd8994: duty=119; 15'd8995: duty=116; 15'd8996: duty=118; 15'd8997: duty=127; 15'd8998: duty=122; 15'd8999: duty=128;
15'd9000: duty=124; 15'd9001: duty=129; 15'd9002: duty=134; 15'd9003: duty=130; 15'd9004: duty=127; 15'd9005: duty=129; 15'd9006: duty=133; 15'd9007: duty=137;
15'd9008: duty=133; 15'd9009: duty=129; 15'd9010: duty=133; 15'd9011: duty=129; 15'd9012: duty=131; 15'd9013: duty=131; 15'd9014: duty=130; 15'd9015: duty=131;
15'd9016: duty=134; 15'd9017: duty=133; 15'd9018: duty=136; 15'd9019: duty=131; 15'd9020: duty=136; 15'd9021: duty=140; 15'd9022: duty=140; 15'd9023: duty=142;
15'd9024: duty=140; 15'd9025: duty=140; 15'd9026: duty=137; 15'd9027: duty=142; 15'd9028: duty=140; 15'd9029: duty=142; 15'd9030: duty=139; 15'd9031: duty=143;
15'd9032: duty=142; 15'd9033: duty=139; 15'd9034: duty=143; 15'd9035: duty=136; 15'd9036: duty=128; 15'd9037: duty=119; 15'd9038: duty=121; 15'd9039: duty=119;
15'd9040: duty=118; 15'd9041: duty=121; 15'd9042: duty=125; 15'd9043: duty=129; 15'd9044: duty=139; 15'd9045: duty=140; 15'd9046: duty=130; 15'd9047: duty=128;
15'd9048: duty=128; 15'd9049: duty=131; 15'd9050: duty=135; 15'd9051: duty=127; 15'd9052: duty=126; 15'd9053: duty=124; 15'd9054: duty=113; 15'd9055: duty=121;
15'd9056: duty=109; 15'd9057: duty=104; 15'd9058: duty=115; 15'd9059: duty=119; 15'd9060: duty=120; 15'd9061: duty=119; 15'd9062: duty=123; 15'd9063: duty=124;
15'd9064: duty=139; 15'd9065: duty=135; 15'd9066: duty=139; 15'd9067: duty=142; 15'd9068: duty=133; 15'd9069: duty=138; 15'd9070: duty=121; 15'd9071: duty=125;
15'd9072: duty=127; 15'd9073: duty=128; 15'd9074: duty=136; 15'd9075: duty=132; 15'd9076: duty=134; 15'd9077: duty=130; 15'd9078: duty=134; 15'd9079: duty=138;
15'd9080: duty=144; 15'd9081: duty=143; 15'd9082: duty=139; 15'd9083: duty=137; 15'd9084: duty=135; 15'd9085: duty=143; 15'd9086: duty=134; 15'd9087: duty=135;
15'd9088: duty=141; 15'd9089: duty=136; 15'd9090: duty=148; 15'd9091: duty=143; 15'd9092: duty=139; 15'd9093: duty=136; 15'd9094: duty=139; 15'd9095: duty=140;
15'd9096: duty=137; 15'd9097: duty=145; 15'd9098: duty=138; 15'd9099: duty=137; 15'd9100: duty=140; 15'd9101: duty=138; 15'd9102: duty=137; 15'd9103: duty=134;
15'd9104: duty=128; 15'd9105: duty=121; 15'd9106: duty=121; 15'd9107: duty=114; 15'd9108: duty=121; 15'd9109: duty=116; 15'd9110: duty=110; 15'd9111: duty=129;
15'd9112: duty=121; 15'd9113: duty=121; 15'd9114: duty=121; 15'd9115: duty=115; 15'd9116: duty=125; 15'd9117: duty=127; 15'd9118: duty=125; 15'd9119: duty=124;
15'd9120: duty=124; 15'd9121: duty=119; 15'd9122: duty=115; 15'd9123: duty=115; 15'd9124: duty=115; 15'd9125: duty=121; 15'd9126: duty=119; 15'd9127: duty=126;
15'd9128: duty=125; 15'd9129: duty=128; 15'd9130: duty=128; 15'd9131: duty=130; 15'd9132: duty=129; 15'd9133: duty=123; 15'd9134: duty=125; 15'd9135: duty=124;
15'd9136: duty=125; 15'd9137: duty=131; 15'd9138: duty=131; 15'd9139: duty=131; 15'd9140: duty=139; 15'd9141: duty=134; 15'd9142: duty=136; 15'd9143: duty=140;
15'd9144: duty=142; 15'd9145: duty=146; 15'd9146: duty=149; 15'd9147: duty=146; 15'd9148: duty=152; 15'd9149: duty=142; 15'd9150: duty=135; 15'd9151: duty=145;
15'd9152: duty=137; 15'd9153: duty=140; 15'd9154: duty=143; 15'd9155: duty=142; 15'd9156: duty=148; 15'd9157: duty=142; 15'd9158: duty=142; 15'd9159: duty=137;
15'd9160: duty=134; 15'd9161: duty=147; 15'd9162: duty=140; 15'd9163: duty=140; 15'd9164: duty=140; 15'd9165: duty=131; 15'd9166: duty=129; 15'd9167: duty=131;
15'd9168: duty=131; 15'd9169: duty=128; 15'd9170: duty=133; 15'd9171: duty=128; 15'd9172: duty=135; 15'd9173: duty=137; 15'd9174: duty=134; 15'd9175: duty=143;
15'd9176: duty=134; 15'd9177: duty=130; 15'd9178: duty=124; 15'd9179: duty=118; 15'd9180: duty=119; 15'd9181: duty=112; 15'd9182: duty=102; 15'd9183: duty=97;
15'd9184: duty=105; 15'd9185: duty=110; 15'd9186: duty=110; 15'd9187: duty=113; 15'd9188: duty=111; 15'd9189: duty=121; 15'd9190: duty=126; 15'd9191: duty=117;
15'd9192: duty=125; 15'd9193: duty=126; 15'd9194: duty=125; 15'd9195: duty=127; 15'd9196: duty=114; 15'd9197: duty=117; 15'd9198: duty=122; 15'd9199: duty=126;
15'd9200: duty=135; 15'd9201: duty=125; 15'd9202: duty=125; 15'd9203: duty=130; 15'd9204: duty=130; 15'd9205: duty=126; 15'd9206: duty=133; 15'd9207: duty=135;
15'd9208: duty=129; 15'd9209: duty=135; 15'd9210: duty=138; 15'd9211: duty=143; 15'd9212: duty=147; 15'd9213: duty=152; 15'd9214: duty=158; 15'd9215: duty=152;
15'd9216: duty=144; 15'd9217: duty=146; 15'd9218: duty=141; 15'd9219: duty=136; 15'd9220: duty=138; 15'd9221: duty=135; 15'd9222: duty=137; 15'd9223: duty=133;
15'd9224: duty=128; 15'd9225: duty=135; 15'd9226: duty=138; 15'd9227: duty=146; 15'd9228: duty=132; 15'd9229: duty=124; 15'd9230: duty=135; 15'd9231: duty=136;
15'd9232: duty=135; 15'd9233: duty=141; 15'd9234: duty=143; 15'd9235: duty=130; 15'd9236: duty=138; 15'd9237: duty=141; 15'd9238: duty=142; 15'd9239: duty=136;
15'd9240: duty=129; 15'd9241: duty=135; 15'd9242: duty=127; 15'd9243: duty=131; 15'd9244: duty=122; 15'd9245: duty=115; 15'd9246: duty=119; 15'd9247: duty=117;
15'd9248: duty=112; 15'd9249: duty=113; 15'd9250: duty=125; 15'd9251: duty=118; 15'd9252: duty=114; 15'd9253: duty=116; 15'd9254: duty=110; 15'd9255: duty=116;
15'd9256: duty=122; 15'd9257: duty=127; 15'd9258: duty=128; 15'd9259: duty=128; 15'd9260: duty=121; 15'd9261: duty=116; 15'd9262: duty=118; 15'd9263: duty=116;
15'd9264: duty=128; 15'd9265: duty=124; 15'd9266: duty=124; 15'd9267: duty=128; 15'd9268: duty=122; 15'd9269: duty=129; 15'd9270: duty=127; 15'd9271: duty=128;
15'd9272: duty=133; 15'd9273: duty=125; 15'd9274: duty=126; 15'd9275: duty=128; 15'd9276: duty=136; 15'd9277: duty=142; 15'd9278: duty=147; 15'd9279: duty=151;
15'd9280: duty=154; 15'd9281: duty=157; 15'd9282: duty=145; 15'd9283: duty=140; 15'd9284: duty=143; 15'd9285: duty=150; 15'd9286: duty=145; 15'd9287: duty=151;
15'd9288: duty=142; 15'd9289: duty=137; 15'd9290: duty=125; 15'd9291: duty=127; 15'd9292: duty=132; 15'd9293: duty=133; 15'd9294: duty=135; 15'd9295: duty=126;
15'd9296: duty=135; 15'd9297: duty=134; 15'd9298: duty=142; 15'd9299: duty=150; 15'd9300: duty=148; 15'd9301: duty=134; 15'd9302: duty=129; 15'd9303: duty=127;
15'd9304: duty=134; 15'd9305: duty=144; 15'd9306: duty=151; 15'd9307: duty=147; 15'd9308: duty=130; 15'd9309: duty=118; 15'd9310: duty=114; 15'd9311: duty=112;
15'd9312: duty=122; 15'd9313: duty=120; 15'd9314: duty=121; 15'd9315: duty=124; 15'd9316: duty=125; 15'd9317: duty=110; 15'd9318: duty=118; 15'd9319: duty=130;
15'd9320: duty=122; 15'd9321: duty=130; 15'd9322: duty=124; 15'd9323: duty=128; 15'd9324: duty=119; 15'd9325: duty=122; 15'd9326: duty=122; 15'd9327: duty=121;
15'd9328: duty=115; 15'd9329: duty=116; 15'd9330: duty=113; 15'd9331: duty=113; 15'd9332: duty=131; 15'd9333: duty=126; 15'd9334: duty=128; 15'd9335: duty=134;
15'd9336: duty=134; 15'd9337: duty=142; 15'd9338: duty=133; 15'd9339: duty=128; 15'd9340: duty=140; 15'd9341: duty=139; 15'd9342: duty=140; 15'd9343: duty=143;
15'd9344: duty=144; 15'd9345: duty=145; 15'd9346: duty=137; 15'd9347: duty=131; 15'd9348: duty=131; 15'd9349: duty=131; 15'd9350: duty=136; 15'd9351: duty=128;
15'd9352: duty=125; 15'd9353: duty=125; 15'd9354: duty=126; 15'd9355: duty=136; 15'd9356: duty=140; 15'd9357: duty=137; 15'd9358: duty=137; 15'd9359: duty=133;
15'd9360: duty=133; 15'd9361: duty=131; 15'd9362: duty=134; 15'd9363: duty=123; 15'd9364: duty=126; 15'd9365: duty=131; 15'd9366: duty=127; 15'd9367: duty=137;
15'd9368: duty=134; 15'd9369: duty=128; 15'd9370: duty=126; 15'd9371: duty=128; 15'd9372: duty=121; 15'd9373: duty=121; 15'd9374: duty=122; 15'd9375: duty=123;
15'd9376: duty=127; 15'd9377: duty=118; 15'd9378: duty=115; 15'd9379: duty=123; 15'd9380: duty=132; 15'd9381: duty=144; 15'd9382: duty=132; 15'd9383: duty=144;
15'd9384: duty=137; 15'd9385: duty=126; 15'd9386: duty=134; 15'd9387: duty=135; 15'd9388: duty=134; 15'd9389: duty=134; 15'd9390: duty=139; 15'd9391: duty=135;
15'd9392: duty=141; 15'd9393: duty=128; 15'd9394: duty=116; 15'd9395: duty=128; 15'd9396: duty=129; 15'd9397: duty=136; 15'd9398: duty=135; 15'd9399: duty=123;
15'd9400: duty=123; 15'd9401: duty=133; 15'd9402: duty=141; 15'd9403: duty=141; 15'd9404: duty=140; 15'd9405: duty=133; 15'd9406: duty=145; 15'd9407: duty=138;
15'd9408: duty=138; 15'd9409: duty=138; 15'd9410: duty=141; 15'd9411: duty=136; 15'd9412: duty=134; 15'd9413: duty=123; 15'd9414: duty=116; 15'd9415: duty=130;
15'd9416: duty=138; 15'd9417: duty=141; 15'd9418: duty=135; 15'd9419: duty=130; 15'd9420: duty=138; 15'd9421: duty=142; 15'd9422: duty=137; 15'd9423: duty=127;
15'd9424: duty=124; 15'd9425: duty=120; 15'd9426: duty=124; 15'd9427: duty=126; 15'd9428: duty=114; 15'd9429: duty=131; 15'd9430: duty=121; 15'd9431: duty=134;
15'd9432: duty=131; 15'd9433: duty=131; 15'd9434: duty=129; 15'd9435: duty=123; 15'd9436: duty=121; 15'd9437: duty=115; 15'd9438: duty=110; 15'd9439: duty=107;
15'd9440: duty=113; 15'd9441: duty=106; 15'd9442: duty=121; 15'd9443: duty=123; 15'd9444: duty=124; 15'd9445: duty=127; 15'd9446: duty=128; 15'd9447: duty=127;
15'd9448: duty=134; 15'd9449: duty=142; 15'd9450: duty=151; 15'd9451: duty=147; 15'd9452: duty=140; 15'd9453: duty=140; 15'd9454: duty=131; 15'd9455: duty=127;
15'd9456: duty=131; 15'd9457: duty=129; 15'd9458: duty=140; 15'd9459: duty=136; 15'd9460: duty=133; 15'd9461: duty=136; 15'd9462: duty=133; 15'd9463: duty=150;
15'd9464: duty=137; 15'd9465: duty=137; 15'd9466: duty=127; 15'd9467: duty=134; 15'd9468: duty=137; 15'd9469: duty=136; 15'd9470: duty=156; 15'd9471: duty=137;
15'd9472: duty=139; 15'd9473: duty=128; 15'd9474: duty=123; 15'd9475: duty=132; 15'd9476: duty=128; 15'd9477: duty=134; 15'd9478: duty=130; 15'd9479: duty=133;
15'd9480: duty=134; 15'd9481: duty=137; 15'd9482: duty=126; 15'd9483: duty=125; 15'd9484: duty=145; 15'd9485: duty=127; 15'd9486: duty=115; 15'd9487: duty=122;
15'd9488: duty=119; 15'd9489: duty=127; 15'd9490: duty=127; 15'd9491: duty=122; 15'd9492: duty=131; 15'd9493: duty=135; 15'd9494: duty=153; 15'd9495: duty=145;
15'd9496: duty=138; 15'd9497: duty=139; 15'd9498: duty=136; 15'd9499: duty=137; 15'd9500: duty=130; 15'd9501: duty=128; 15'd9502: duty=116; 15'd9503: duty=110;
15'd9504: duty=119; 15'd9505: duty=110; 15'd9506: duty=104; 15'd9507: duty=118; 15'd9508: duty=128; 15'd9509: duty=127; 15'd9510: duty=121; 15'd9511: duty=124;
15'd9512: duty=118; 15'd9513: duty=129; 15'd9514: duty=134; 15'd9515: duty=137; 15'd9516: duty=127; 15'd9517: duty=127; 15'd9518: duty=133; 15'd9519: duty=124;
15'd9520: duty=128; 15'd9521: duty=134; 15'd9522: duty=137; 15'd9523: duty=136; 15'd9524: duty=142; 15'd9525: duty=134; 15'd9526: duty=146; 15'd9527: duty=125;
15'd9528: duty=127; 15'd9529: duty=140; 15'd9530: duty=139; 15'd9531: duty=139; 15'd9532: duty=131; 15'd9533: duty=140; 15'd9534: duty=140; 15'd9535: duty=145;
15'd9536: duty=131; 15'd9537: duty=142; 15'd9538: duty=134; 15'd9539: duty=133; 15'd9540: duty=140; 15'd9541: duty=133; 15'd9542: duty=148; 15'd9543: duty=137;
15'd9544: duty=143; 15'd9545: duty=134; 15'd9546: duty=126; 15'd9547: duty=128; 15'd9548: duty=123; 15'd9549: duty=124; 15'd9550: duty=104; 15'd9551: duty=113;
15'd9552: duty=124; 15'd9553: duty=119; 15'd9554: duty=121; 15'd9555: duty=128; 15'd9556: duty=139; 15'd9557: duty=135; 15'd9558: duty=148; 15'd9559: duty=136;
15'd9560: duty=127; 15'd9561: duty=134; 15'd9562: duty=131; 15'd9563: duty=142; 15'd9564: duty=131; 15'd9565: duty=128; 15'd9566: duty=127; 15'd9567: duty=128;
15'd9568: duty=121; 15'd9569: duty=110; 15'd9570: duty=113; 15'd9571: duty=106; 15'd9572: duty=112; 15'd9573: duty=116; 15'd9574: duty=128; 15'd9575: duty=124;
15'd9576: duty=122; 15'd9577: duty=145; 15'd9578: duty=143; 15'd9579: duty=150; 15'd9580: duty=143; 15'd9581: duty=145; 15'd9582: duty=150; 15'd9583: duty=147;
15'd9584: duty=148; 15'd9585: duty=133; 15'd9586: duty=124; 15'd9587: duty=127; 15'd9588: duty=130; 15'd9589: duty=133; 15'd9590: duty=137; 15'd9591: duty=137;
15'd9592: duty=142; 15'd9593: duty=148; 15'd9594: duty=150; 15'd9595: duty=146; 15'd9596: duty=142; 15'd9597: duty=138; 15'd9598: duty=147; 15'd9599: duty=140;
15'd9600: duty=148; 15'd9601: duty=154; 15'd9602: duty=142; 15'd9603: duty=143; 15'd9604: duty=121; 15'd9605: duty=124; 15'd9606: duty=123; 15'd9607: duty=124;
15'd9608: duty=134; 15'd9609: duty=119; 15'd9610: duty=130; 15'd9611: duty=120; 15'd9612: duty=120; 15'd9613: duty=117; 15'd9614: duty=110; 15'd9615: duty=122;
15'd9616: duty=124; 15'd9617: duty=124; 15'd9618: duty=109; 15'd9619: duty=113; 15'd9620: duty=112; 15'd9621: duty=117; 15'd9622: duty=127; 15'd9623: duty=118;
15'd9624: duty=128; 15'd9625: duty=127; 15'd9626: duty=121; 15'd9627: duty=121; 15'd9628: duty=119; 15'd9629: duty=121; 15'd9630: duty=124; 15'd9631: duty=123;
15'd9632: duty=109; 15'd9633: duty=109; 15'd9634: duty=115; 15'd9635: duty=118; 15'd9636: duty=127; 15'd9637: duty=123; 15'd9638: duty=131; 15'd9639: duty=133;
15'd9640: duty=114; 15'd9641: duty=123; 15'd9642: duty=120; 15'd9643: duty=124; 15'd9644: duty=132; 15'd9645: duty=145; 15'd9646: duty=139; 15'd9647: duty=141;
15'd9648: duty=149; 15'd9649: duty=151; 15'd9650: duty=152; 15'd9651: duty=130; 15'd9652: duty=127; 15'd9653: duty=130; 15'd9654: duty=141; 15'd9655: duty=136;
15'd9656: duty=146; 15'd9657: duty=150; 15'd9658: duty=156; 15'd9659: duty=151; 15'd9660: duty=150; 15'd9661: duty=163; 15'd9662: duty=159; 15'd9663: duty=151;
15'd9664: duty=151; 15'd9665: duty=145; 15'd9666: duty=139; 15'd9667: duty=137; 15'd9668: duty=122; 15'd9669: duty=148; 15'd9670: duty=147; 15'd9671: duty=138;
15'd9672: duty=138; 15'd9673: duty=129; 15'd9674: duty=132; 15'd9675: duty=132; 15'd9676: duty=135; 15'd9677: duty=143; 15'd9678: duty=133; 15'd9679: duty=129;
15'd9680: duty=131; 15'd9681: duty=122; 15'd9682: duty=126; 15'd9683: duty=114; 15'd9684: duty=109; 15'd9685: duty=110; 15'd9686: duty=108; 15'd9687: duty=105;
15'd9688: duty=107; 15'd9689: duty=125; 15'd9690: duty=130; 15'd9691: duty=125; 15'd9692: duty=127; 15'd9693: duty=130; 15'd9694: duty=138; 15'd9695: duty=143;
15'd9696: duty=147; 15'd9697: duty=138; 15'd9698: duty=120; 15'd9699: duty=122; 15'd9700: duty=114; 15'd9701: duty=100; 15'd9702: duty=95; 15'd9703: duty=105;
15'd9704: duty=114; 15'd9705: duty=111; 15'd9706: duty=114; 15'd9707: duty=110; 15'd9708: duty=127; 15'd9709: duty=128; 15'd9710: duty=127; 15'd9711: duty=130;
15'd9712: duty=123; 15'd9713: duty=141; 15'd9714: duty=144; 15'd9715: duty=146; 15'd9716: duty=147; 15'd9717: duty=142; 15'd9718: duty=136; 15'd9719: duty=149;
15'd9720: duty=145; 15'd9721: duty=142; 15'd9722: duty=144; 15'd9723: duty=136; 15'd9724: duty=149; 15'd9725: duty=136; 15'd9726: duty=130; 15'd9727: duty=140;
15'd9728: duty=153; 15'd9729: duty=149; 15'd9730: duty=154; 15'd9731: duty=153; 15'd9732: duty=142; 15'd9733: duty=146; 15'd9734: duty=139; 15'd9735: duty=137;
15'd9736: duty=127; 15'd9737: duty=134; 15'd9738: duty=127; 15'd9739: duty=99; 15'd9740: duty=107; 15'd9741: duty=119; 15'd9742: duty=110; 15'd9743: duty=115;
15'd9744: duty=118; 15'd9745: duty=127; 15'd9746: duty=125; 15'd9747: duty=125; 15'd9748: duty=125; 15'd9749: duty=121; 15'd9750: duty=126; 15'd9751: duty=131;
15'd9752: duty=134; 15'd9753: duty=139; 15'd9754: duty=131; 15'd9755: duty=116; 15'd9756: duty=124; 15'd9757: duty=126; 15'd9758: duty=119; 15'd9759: duty=108;
15'd9760: duty=115; 15'd9761: duty=124; 15'd9762: duty=144; 15'd9763: duty=139; 15'd9764: duty=132; 15'd9765: duty=122; 15'd9766: duty=115; 15'd9767: duty=122;
15'd9768: duty=117; 15'd9769: duty=119; 15'd9770: duty=124; 15'd9771: duty=140; 15'd9772: duty=148; 15'd9773: duty=133; 15'd9774: duty=133; 15'd9775: duty=128;
15'd9776: duty=127; 15'd9777: duty=140; 15'd9778: duty=132; 15'd9779: duty=136; 15'd9780: duty=133; 15'd9781: duty=126; 15'd9782: duty=135; 15'd9783: duty=141;
15'd9784: duty=141; 15'd9785: duty=155; 15'd9786: duty=147; 15'd9787: duty=146; 15'd9788: duty=149; 15'd9789: duty=144; 15'd9790: duty=144; 15'd9791: duty=163;
15'd9792: duty=159; 15'd9793: duty=154; 15'd9794: duty=142; 15'd9795: duty=128; 15'd9796: duty=126; 15'd9797: duty=123; 15'd9798: duty=142; 15'd9799: duty=138;
15'd9800: duty=136; 15'd9801: duty=127; 15'd9802: duty=138; 15'd9803: duty=129; 15'd9804: duty=153; 15'd9805: duty=140; 15'd9806: duty=150; 15'd9807: duty=148;
15'd9808: duty=121; 15'd9809: duty=137; 15'd9810: duty=123; 15'd9811: duty=127; 15'd9812: duty=110; 15'd9813: duty=121; 15'd9814: duty=110; 15'd9815: duty=101;
15'd9816: duty=110; 15'd9817: duty=107; 15'd9818: duty=104; 15'd9819: duty=121; 15'd9820: duty=133; 15'd9821: duty=127; 15'd9822: duty=119; 15'd9823: duty=124;
15'd9824: duty=121; 15'd9825: duty=128; 15'd9826: duty=128; 15'd9827: duty=113; 15'd9828: duty=104; 15'd9829: duty=112; 15'd9830: duty=119; 15'd9831: duty=111;
15'd9832: duty=122; 15'd9833: duty=107; 15'd9834: duty=110; 15'd9835: duty=109; 15'd9836: duty=113; 15'd9837: duty=109; 15'd9838: duty=114; 15'd9839: duty=130;
15'd9840: duty=134; 15'd9841: duty=129; 15'd9842: duty=138; 15'd9843: duty=139; 15'd9844: duty=127; 15'd9845: duty=145; 15'd9846: duty=146; 15'd9847: duty=139;
15'd9848: duty=140; 15'd9849: duty=140; 15'd9850: duty=142; 15'd9851: duty=152; 15'd9852: duty=146; 15'd9853: duty=151; 15'd9854: duty=156; 15'd9855: duty=159;
15'd9856: duty=155; 15'd9857: duty=159; 15'd9858: duty=155; 15'd9859: duty=153; 15'd9860: duty=146; 15'd9861: duty=139; 15'd9862: duty=140; 15'd9863: duty=133;
15'd9864: duty=147; 15'd9865: duty=154; 15'd9866: duty=146; 15'd9867: duty=153; 15'd9868: duty=154; 15'd9869: duty=150; 15'd9870: duty=141; 15'd9871: duty=128;
15'd9872: duty=138; 15'd9873: duty=123; 15'd9874: duty=132; 15'd9875: duty=124; 15'd9876: duty=128; 15'd9877: duty=124; 15'd9878: duty=121; 15'd9879: duty=119;
15'd9880: duty=119; 15'd9881: duty=126; 15'd9882: duty=125; 15'd9883: duty=126; 15'd9884: duty=117; 15'd9885: duty=113; 15'd9886: duty=102; 15'd9887: duty=107;
15'd9888: duty=101; 15'd9889: duty=109; 15'd9890: duty=107; 15'd9891: duty=96; 15'd9892: duty=95; 15'd9893: duty=105; 15'd9894: duty=106; 15'd9895: duty=110;
15'd9896: duty=107; 15'd9897: duty=113; 15'd9898: duty=113; 15'd9899: duty=118; 15'd9900: duty=122; 15'd9901: duty=125; 15'd9902: duty=124; 15'd9903: duty=130;
15'd9904: duty=121; 15'd9905: duty=127; 15'd9906: duty=133; 15'd9907: duty=121; 15'd9908: duty=128; 15'd9909: duty=136; 15'd9910: duty=136; 15'd9911: duty=140;
15'd9912: duty=145; 15'd9913: duty=130; 15'd9914: duty=136; 15'd9915: duty=137; 15'd9916: duty=139; 15'd9917: duty=134; 15'd9918: duty=137; 15'd9919: duty=140;
15'd9920: duty=150; 15'd9921: duty=149; 15'd9922: duty=155; 15'd9923: duty=149; 15'd9924: duty=159; 15'd9925: duty=159; 15'd9926: duty=152; 15'd9927: duty=151;
15'd9928: duty=149; 15'd9929: duty=140; 15'd9930: duty=140; 15'd9931: duty=143; 15'd9932: duty=140; 15'd9933: duty=145; 15'd9934: duty=149; 15'd9935: duty=152;
15'd9936: duty=147; 15'd9937: duty=159; 15'd9938: duty=140; 15'd9939: duty=138; 15'd9940: duty=130; 15'd9941: duty=134; 15'd9942: duty=136; 15'd9943: duty=136;
15'd9944: duty=140; 15'd9945: duty=134; 15'd9946: duty=121; 15'd9947: duty=128; 15'd9948: duty=128; 15'd9949: duty=119; 15'd9950: duty=124; 15'd9951: duty=119;
15'd9952: duty=126; 15'd9953: duty=129; 15'd9954: duty=133; 15'd9955: duty=113; 15'd9956: duty=109; 15'd9957: duty=119; 15'd9958: duty=111; 15'd9959: duty=107;
15'd9960: duty=96; 15'd9961: duty=104; 15'd9962: duty=124; 15'd9963: duty=128; 15'd9964: duty=119; 15'd9965: duty=127; 15'd9966: duty=118; 15'd9967: duty=111;
15'd9968: duty=109; 15'd9969: duty=103; 15'd9970: duty=106; 15'd9971: duty=111; 15'd9972: duty=116; 15'd9973: duty=110; 15'd9974: duty=116; 15'd9975: duty=126;
15'd9976: duty=128; 15'd9977: duty=119; 15'd9978: duty=126; 15'd9979: duty=138; 15'd9980: duty=134; 15'd9981: duty=140; 15'd9982: duty=144; 15'd9983: duty=142;
15'd9984: duty=141; 15'd9985: duty=134; 15'd9986: duty=139; 15'd9987: duty=145; 15'd9988: duty=147; 15'd9989: duty=153; 15'd9990: duty=153; 15'd9991: duty=138;
15'd9992: duty=144; 15'd9993: duty=150; 15'd9994: duty=138; 15'd9995: duty=141; 15'd9996: duty=138; 15'd9997: duty=142; 15'd9998: duty=147; 15'd9999: duty=150;
15'd10000: duty=151; 15'd10001: duty=150; 15'd10002: duty=148; 15'd10003: duty=136; 15'd10004: duty=136; 15'd10005: duty=145; 15'd10006: duty=151; 15'd10007: duty=146;
15'd10008: duty=145; 15'd10009: duty=129; 15'd10010: duty=126; 15'd10011: duty=131; 15'd10012: duty=131; 15'd10013: duty=126; 15'd10014: duty=127; 15'd10015: duty=129;
15'd10016: duty=119; 15'd10017: duty=121; 15'd10018: duty=121; 15'd10019: duty=127; 15'd10020: duty=119; 15'd10021: duty=115; 15'd10022: duty=116; 15'd10023: duty=129;
15'd10024: duty=119; 15'd10025: duty=116; 15'd10026: duty=116; 15'd10027: duty=118; 15'd10028: duty=124; 15'd10029: duty=128; 15'd10030: duty=111; 15'd10031: duty=101;
15'd10032: duty=110; 15'd10033: duty=114; 15'd10034: duty=122; 15'd10035: duty=121; 15'd10036: duty=124; 15'd10037: duty=130; 15'd10038: duty=133; 15'd10039: duty=131;
15'd10040: duty=129; 15'd10041: duty=135; 15'd10042: duty=137; 15'd10043: duty=125; 15'd10044: duty=128; 15'd10045: duty=125; 15'd10046: duty=118; 15'd10047: duty=125;
15'd10048: duty=129; 15'd10049: duty=124; 15'd10050: duty=144; 15'd10051: duty=140; 15'd10052: duty=137; 15'd10053: duty=141; 15'd10054: duty=148; 15'd10055: duty=149;
15'd10056: duty=148; 15'd10057: duty=146; 15'd10058: duty=140; 15'd10059: duty=143; 15'd10060: duty=151; 15'd10061: duty=143; 15'd10062: duty=129; 15'd10063: duty=133;
15'd10064: duty=131; 15'd10065: duty=129; 15'd10066: duty=144; 15'd10067: duty=153; 15'd10068: duty=147; 15'd10069: duty=151; 15'd10070: duty=148; 15'd10071: duty=142;
15'd10072: duty=131; 15'd10073: duty=133; 15'd10074: duty=147; 15'd10075: duty=139; 15'd10076: duty=133; 15'd10077: duty=127; 15'd10078: duty=128; 15'd10079: duty=141;
15'd10080: duty=122; 15'd10081: duty=118; 15'd10082: duty=115; 15'd10083: duty=123; 15'd10084: duty=127; 15'd10085: duty=127; 15'd10086: duty=132; 15'd10087: duty=118;
15'd10088: duty=119; 15'd10089: duty=121; 15'd10090: duty=122; 15'd10091: duty=124; 15'd10092: duty=110; 15'd10093: duty=126; 15'd10094: duty=111; 15'd10095: duty=111;
15'd10096: duty=108; 15'd10097: duty=117; 15'd10098: duty=140; 15'd10099: duty=120; 15'd10100: duty=122; 15'd10101: duty=122; 15'd10102: duty=119; 15'd10103: duty=107;
15'd10104: duty=114; 15'd10105: duty=107; 15'd10106: duty=111; 15'd10107: duty=121; 15'd10108: duty=122; 15'd10109: duty=119; 15'd10110: duty=119; 15'd10111: duty=126;
15'd10112: duty=119; 15'd10113: duty=121; 15'd10114: duty=132; 15'd10115: duty=125; 15'd10116: duty=141; 15'd10117: duty=142; 15'd10118: duty=137; 15'd10119: duty=141;
15'd10120: duty=141; 15'd10121: duty=145; 15'd10122: duty=147; 15'd10123: duty=134; 15'd10124: duty=130; 15'd10125: duty=142; 15'd10126: duty=139; 15'd10127: duty=146;
15'd10128: duty=141; 15'd10129: duty=131; 15'd10130: duty=141; 15'd10131: duty=153; 15'd10132: duty=145; 15'd10133: duty=148; 15'd10134: duty=144; 15'd10135: duty=144;
15'd10136: duty=140; 15'd10137: duty=150; 15'd10138: duty=152; 15'd10139: duty=152; 15'd10140: duty=147; 15'd10141: duty=145; 15'd10142: duty=146; 15'd10143: duty=143;
15'd10144: duty=136; 15'd10145: duty=134; 15'd10146: duty=139; 15'd10147: duty=134; 15'd10148: duty=128; 15'd10149: duty=128; 15'd10150: duty=122; 15'd10151: duty=121;
15'd10152: duty=122; 15'd10153: duty=115; 15'd10154: duty=126; 15'd10155: duty=121; 15'd10156: duty=129; 15'd10157: duty=124; 15'd10158: duty=127; 15'd10159: duty=122;
15'd10160: duty=123; 15'd10161: duty=121; 15'd10162: duty=122; 15'd10163: duty=128; 15'd10164: duty=115; 15'd10165: duty=120; 15'd10166: duty=114; 15'd10167: duty=102;
15'd10168: duty=116; 15'd10169: duty=110; 15'd10170: duty=101; 15'd10171: duty=112; 15'd10172: duty=112; 15'd10173: duty=121; 15'd10174: duty=121; 15'd10175: duty=134;
15'd10176: duty=133; 15'd10177: duty=127; 15'd10178: duty=140; 15'd10179: duty=131; 15'd10180: duty=135; 15'd10181: duty=142; 15'd10182: duty=132; 15'd10183: duty=131;
15'd10184: duty=116; 15'd10185: duty=127; 15'd10186: duty=126; 15'd10187: duty=120; 15'd10188: duty=127; 15'd10189: duty=130; 15'd10190: duty=131; 15'd10191: duty=137;
15'd10192: duty=142; 15'd10193: duty=150; 15'd10194: duty=151; 15'd10195: duty=136; 15'd10196: duty=142; 15'd10197: duty=137; 15'd10198: duty=131; 15'd10199: duty=128;
15'd10200: duty=133; 15'd10201: duty=136; 15'd10202: duty=144; 15'd10203: duty=144; 15'd10204: duty=146; 15'd10205: duty=143; 15'd10206: duty=137; 15'd10207: duty=139;
15'd10208: duty=142; 15'd10209: duty=148; 15'd10210: duty=148; 15'd10211: duty=151; 15'd10212: duty=144; 15'd10213: duty=141; 15'd10214: duty=139; 15'd10215: duty=136;
15'd10216: duty=132; 15'd10217: duty=120; 15'd10218: duty=125; 15'd10219: duty=128; 15'd10220: duty=129; 15'd10221: duty=115; 15'd10222: duty=122; 15'd10223: duty=128;
15'd10224: duty=132; 15'd10225: duty=151; 15'd10226: duty=139; 15'd10227: duty=145; 15'd10228: duty=122; 15'd10229: duty=98; 15'd10230: duty=107; 15'd10231: duty=113;
15'd10232: duty=121; 15'd10233: duty=128; 15'd10234: duty=122; 15'd10235: duty=128; 15'd10236: duty=125; 15'd10237: duty=124; 15'd10238: duty=114; 15'd10239: duty=112;
15'd10240: duty=118; 15'd10241: duty=125; 15'd10242: duty=128; 15'd10243: duty=133; 15'd10244: duty=137; 15'd10245: duty=127; 15'd10246: duty=133; 15'd10247: duty=124;
15'd10248: duty=116; 15'd10249: duty=113; 15'd10250: duty=112; 15'd10251: duty=118; 15'd10252: duty=129; 15'd10253: duty=128; 15'd10254: duty=133; 15'd10255: duty=127;
15'd10256: duty=121; 15'd10257: duty=121; 15'd10258: duty=117; 15'd10259: duty=133; 15'd10260: duty=144; 15'd10261: duty=146; 15'd10262: duty=147; 15'd10263: duty=153;
15'd10264: duty=153; 15'd10265: duty=154; 15'd10266: duty=150; 15'd10267: duty=134; 15'd10268: duty=133; 15'd10269: duty=127; 15'd10270: duty=127; 15'd10271: duty=143;
15'd10272: duty=148; 15'd10273: duty=154; 15'd10274: duty=156; 15'd10275: duty=158; 15'd10276: duty=154; 15'd10277: duty=147; 15'd10278: duty=145; 15'd10279: duty=142;
15'd10280: duty=141; 15'd10281: duty=136; 15'd10282: duty=141; 15'd10283: duty=144; 15'd10284: duty=131; 15'd10285: duty=127; 15'd10286: duty=122; 15'd10287: duty=118;
15'd10288: duty=116; 15'd10289: duty=112; 15'd10290: duty=125; 15'd10291: duty=135; 15'd10292: duty=125; 15'd10293: duty=122; 15'd10294: duty=119; 15'd10295: duty=104;
15'd10296: duty=109; 15'd10297: duty=107; 15'd10298: duty=103; 15'd10299: duty=109; 15'd10300: duty=120; 15'd10301: duty=118; 15'd10302: duty=119; 15'd10303: duty=127;
15'd10304: duty=125; 15'd10305: duty=114; 15'd10306: duty=117; 15'd10307: duty=119; 15'd10308: duty=116; 15'd10309: duty=136; 15'd10310: duty=122; 15'd10311: duty=126;
15'd10312: duty=124; 15'd10313: duty=119; 15'd10314: duty=134; 15'd10315: duty=129; 15'd10316: duty=132; 15'd10317: duty=144; 15'd10318: duty=145; 15'd10319: duty=139;
15'd10320: duty=142; 15'd10321: duty=145; 15'd10322: duty=143; 15'd10323: duty=138; 15'd10324: duty=136; 15'd10325: duty=128; 15'd10326: duty=124; 15'd10327: duty=128;
15'd10328: duty=128; 15'd10329: duty=126; 15'd10330: duty=124; 15'd10331: duty=127; 15'd10332: duty=138; 15'd10333: duty=145; 15'd10334: duty=149; 15'd10335: duty=148;
15'd10336: duty=144; 15'd10337: duty=145; 15'd10338: duty=148; 15'd10339: duty=144; 15'd10340: duty=145; 15'd10341: duty=143; 15'd10342: duty=144; 15'd10343: duty=137;
15'd10344: duty=135; 15'd10345: duty=148; 15'd10346: duty=144; 15'd10347: duty=143; 15'd10348: duty=131; 15'd10349: duty=126; 15'd10350: duty=131; 15'd10351: duty=138;
15'd10352: duty=141; 15'd10353: duty=130; 15'd10354: duty=123; 15'd10355: duty=130; 15'd10356: duty=123; 15'd10357: duty=126; 15'd10358: duty=133; 15'd10359: duty=122;
15'd10360: duty=126; 15'd10361: duty=119; 15'd10362: duty=124; 15'd10363: duty=119; 15'd10364: duty=109; 15'd10365: duty=110; 15'd10366: duty=117; 15'd10367: duty=134;
15'd10368: duty=130; 15'd10369: duty=110; 15'd10370: duty=117; 15'd10371: duty=118; 15'd10372: duty=116; 15'd10373: duty=127; 15'd10374: duty=127; 15'd10375: duty=129;
15'd10376: duty=121; 15'd10377: duty=122; 15'd10378: duty=115; 15'd10379: duty=127; 15'd10380: duty=133; 15'd10381: duty=110; 15'd10382: duty=113; 15'd10383: duty=134;
15'd10384: duty=132; 15'd10385: duty=121; 15'd10386: duty=124; 15'd10387: duty=130; 15'd10388: duty=130; 15'd10389: duty=136; 15'd10390: duty=137; 15'd10391: duty=125;
15'd10392: duty=135; 15'd10393: duty=134; 15'd10394: duty=133; 15'd10395: duty=150; 15'd10396: duty=144; 15'd10397: duty=129; 15'd10398: duty=127; 15'd10399: duty=132;
15'd10400: duty=136; 15'd10401: duty=140; 15'd10402: duty=151; 15'd10403: duty=142; 15'd10404: duty=139; 15'd10405: duty=147; 15'd10406: duty=144; 15'd10407: duty=144;
15'd10408: duty=139; 15'd10409: duty=137; 15'd10410: duty=139; 15'd10411: duty=140; 15'd10412: duty=139; 15'd10413: duty=146; 15'd10414: duty=145; 15'd10415: duty=143;
15'd10416: duty=142; 15'd10417: duty=128; 15'd10418: duty=138; 15'd10419: duty=144; 15'd10420: duty=145; 15'd10421: duty=148; 15'd10422: duty=136; 15'd10423: duty=137;
15'd10424: duty=133; 15'd10425: duty=125; 15'd10426: duty=127; 15'd10427: duty=131; 15'd10428: duty=124; 15'd10429: duty=116; 15'd10430: duty=126; 15'd10431: duty=132;
15'd10432: duty=110; 15'd10433: duty=116; 15'd10434: duty=123; 15'd10435: duty=119; 15'd10436: duty=109; 15'd10437: duty=108; 15'd10438: duty=115; 15'd10439: duty=114;
15'd10440: duty=116; 15'd10441: duty=109; 15'd10442: duty=118; 15'd10443: duty=118; 15'd10444: duty=109; 15'd10445: duty=102; 15'd10446: duty=105; 15'd10447: duty=107;
15'd10448: duty=121; 15'd10449: duty=113; 15'd10450: duty=118; 15'd10451: duty=131; 15'd10452: duty=133; 15'd10453: duty=143; 15'd10454: duty=143; 15'd10455: duty=148;
15'd10456: duty=140; 15'd10457: duty=133; 15'd10458: duty=130; 15'd10459: duty=125; 15'd10460: duty=125; 15'd10461: duty=131; 15'd10462: duty=131; 15'd10463: duty=143;
15'd10464: duty=153; 15'd10465: duty=148; 15'd10466: duty=150; 15'd10467: duty=149; 15'd10468: duty=148; 15'd10469: duty=141; 15'd10470: duty=134; 15'd10471: duty=130;
15'd10472: duty=127; 15'd10473: duty=126; 15'd10474: duty=131; 15'd10475: duty=135; 15'd10476: duty=133; 15'd10477: duty=130; 15'd10478: duty=127; 15'd10479: duty=135;
15'd10480: duty=145; 15'd10481: duty=136; 15'd10482: duty=132; 15'd10483: duty=139; 15'd10484: duty=141; 15'd10485: duty=145; 15'd10486: duty=144; 15'd10487: duty=147;
15'd10488: duty=140; 15'd10489: duty=145; 15'd10490: duty=143; 15'd10491: duty=151; 15'd10492: duty=145; 15'd10493: duty=136; 15'd10494: duty=132; 15'd10495: duty=129;
15'd10496: duty=143; 15'd10497: duty=128; 15'd10498: duty=128; 15'd10499: duty=122; 15'd10500: duty=125; 15'd10501: duty=108; 15'd10502: duty=105; 15'd10503: duty=104;
15'd10504: duty=111; 15'd10505: duty=127; 15'd10506: duty=114; 15'd10507: duty=122; 15'd10508: duty=138; 15'd10509: duty=131; 15'd10510: duty=120; 15'd10511: duty=122;
15'd10512: duty=126; 15'd10513: duty=128; 15'd10514: duty=126; 15'd10515: duty=120; 15'd10516: duty=114; 15'd10517: duty=127; 15'd10518: duty=117; 15'd10519: duty=110;
15'd10520: duty=111; 15'd10521: duty=110; 15'd10522: duty=107; 15'd10523: duty=113; 15'd10524: duty=115; 15'd10525: duty=116; 15'd10526: duty=122; 15'd10527: duty=122;
15'd10528: duty=121; 15'd10529: duty=121; 15'd10530: duty=124; 15'd10531: duty=129; 15'd10532: duty=136; 15'd10533: duty=136; 15'd10534: duty=139; 15'd10535: duty=147;
15'd10536: duty=149; 15'd10537: duty=150; 15'd10538: duty=142; 15'd10539: duty=140; 15'd10540: duty=143; 15'd10541: duty=128; 15'd10542: duty=131; 15'd10543: duty=143;
15'd10544: duty=142; 15'd10545: duty=135; 15'd10546: duty=150; 15'd10547: duty=152; 15'd10548: duty=148; 15'd10549: duty=157; 15'd10550: duty=147; 15'd10551: duty=143;
15'd10552: duty=142; 15'd10553: duty=141; 15'd10554: duty=145; 15'd10555: duty=151; 15'd10556: duty=148; 15'd10557: duty=151; 15'd10558: duty=138; 15'd10559: duty=140;
15'd10560: duty=149; 15'd10561: duty=141; 15'd10562: duty=143; 15'd10563: duty=129; 15'd10564: duty=141; 15'd10565: duty=133; 15'd10566: duty=126; 15'd10567: duty=136;
15'd10568: duty=123; 15'd10569: duty=129; 15'd10570: duty=127; 15'd10571: duty=130; 15'd10572: duty=132; 15'd10573: duty=135; 15'd10574: duty=130; 15'd10575: duty=120;
15'd10576: duty=121; 15'd10577: duty=113; 15'd10578: duty=117; 15'd10579: duty=114; 15'd10580: duty=112; 15'd10581: duty=112; 15'd10582: duty=104; 15'd10583: duty=105;
15'd10584: duty=108; 15'd10585: duty=111; 15'd10586: duty=106; 15'd10587: duty=125; 15'd10588: duty=116; 15'd10589: duty=111; 15'd10590: duty=127; 15'd10591: duty=125;
15'd10592: duty=123; 15'd10593: duty=117; 15'd10594: duty=117; 15'd10595: duty=122; 15'd10596: duty=126; 15'd10597: duty=126; 15'd10598: duty=114; 15'd10599: duty=120;
15'd10600: duty=135; 15'd10601: duty=122; 15'd10602: duty=133; 15'd10603: duty=146; 15'd10604: duty=139; 15'd10605: duty=135; 15'd10606: duty=148; 15'd10607: duty=149;
15'd10608: duty=149; 15'd10609: duty=154; 15'd10610: duty=149; 15'd10611: duty=145; 15'd10612: duty=137; 15'd10613: duty=134; 15'd10614: duty=142; 15'd10615: duty=141;
15'd10616: duty=136; 15'd10617: duty=137; 15'd10618: duty=129; 15'd10619: duty=134; 15'd10620: duty=141; 15'd10621: duty=141; 15'd10622: duty=134; 15'd10623: duty=146;
15'd10624: duty=150; 15'd10625: duty=156; 15'd10626: duty=155; 15'd10627: duty=144; 15'd10628: duty=134; 15'd10629: duty=136; 15'd10630: duty=140; 15'd10631: duty=138;
15'd10632: duty=141; 15'd10633: duty=139; 15'd10634: duty=142; 15'd10635: duty=139; 15'd10636: duty=132; 15'd10637: duty=121; 15'd10638: duty=124; 15'd10639: duty=120;
15'd10640: duty=123; 15'd10641: duty=119; 15'd10642: duty=129; 15'd10643: duty=134; 15'd10644: duty=126; 15'd10645: duty=114; 15'd10646: duty=110; 15'd10647: duty=117;
15'd10648: duty=119; 15'd10649: duty=117; 15'd10650: duty=118; 15'd10651: duty=125; 15'd10652: duty=120; 15'd10653: duty=135; 15'd10654: duty=130; 15'd10655: duty=125;
15'd10656: duty=118; 15'd10657: duty=111; 15'd10658: duty=107; 15'd10659: duty=110; 15'd10660: duty=106; 15'd10661: duty=108; 15'd10662: duty=118; 15'd10663: duty=114;
15'd10664: duty=107; 15'd10665: duty=107; 15'd10666: duty=115; 15'd10667: duty=115; 15'd10668: duty=121; 15'd10669: duty=124; 15'd10670: duty=131; 15'd10671: duty=130;
15'd10672: duty=133; 15'd10673: duty=128; 15'd10674: duty=133; 15'd10675: duty=136; 15'd10676: duty=133; 15'd10677: duty=131; 15'd10678: duty=130; 15'd10679: duty=143;
15'd10680: duty=136; 15'd10681: duty=131; 15'd10682: duty=139; 15'd10683: duty=145; 15'd10684: duty=150; 15'd10685: duty=147; 15'd10686: duty=147; 15'd10687: duty=143;
15'd10688: duty=147; 15'd10689: duty=154; 15'd10690: duty=147; 15'd10691: duty=148; 15'd10692: duty=136; 15'd10693: duty=143; 15'd10694: duty=144; 15'd10695: duty=140;
15'd10696: duty=142; 15'd10697: duty=149; 15'd10698: duty=145; 15'd10699: duty=148; 15'd10700: duty=146; 15'd10701: duty=140; 15'd10702: duty=145; 15'd10703: duty=143;
15'd10704: duty=141; 15'd10705: duty=150; 15'd10706: duty=144; 15'd10707: duty=130; 15'd10708: duty=139; 15'd10709: duty=132; 15'd10710: duty=130; 15'd10711: duty=126;
15'd10712: duty=127; 15'd10713: duty=128; 15'd10714: duty=132; 15'd10715: duty=138; 15'd10716: duty=137; 15'd10717: duty=129; 15'd10718: duty=129; 15'd10719: duty=126;
15'd10720: duty=127; 15'd10721: duty=121; 15'd10722: duty=104; 15'd10723: duty=103; 15'd10724: duty=107; 15'd10725: duty=112; 15'd10726: duty=114; 15'd10727: duty=123;
15'd10728: duty=122; 15'd10729: duty=115; 15'd10730: duty=119; 15'd10731: duty=118; 15'd10732: duty=113; 15'd10733: duty=114; 15'd10734: duty=104; 15'd10735: duty=108;
15'd10736: duty=107; 15'd10737: duty=109; 15'd10738: duty=111; 15'd10739: duty=104; 15'd10740: duty=103; 15'd10741: duty=111; 15'd10742: duty=117; 15'd10743: duty=118;
15'd10744: duty=127; 15'd10745: duty=133; 15'd10746: duty=123; 15'd10747: duty=118; 15'd10748: duty=119; 15'd10749: duty=124; 15'd10750: duty=131; 15'd10751: duty=133;
15'd10752: duty=131; 15'd10753: duty=134; 15'd10754: duty=148; 15'd10755: duty=143; 15'd10756: duty=150; 15'd10757: duty=145; 15'd10758: duty=147; 15'd10759: duty=151;
15'd10760: duty=155; 15'd10761: duty=163; 15'd10762: duty=152; 15'd10763: duty=147; 15'd10764: duty=150; 15'd10765: duty=152; 15'd10766: duty=147; 15'd10767: duty=154;
15'd10768: duty=150; 15'd10769: duty=151; 15'd10770: duty=146; 15'd10771: duty=146; 15'd10772: duty=148; 15'd10773: duty=151; 15'd10774: duty=161; 15'd10775: duty=155;
15'd10776: duty=151; 15'd10777: duty=152; 15'd10778: duty=151; 15'd10779: duty=146; 15'd10780: duty=144; 15'd10781: duty=135; 15'd10782: duty=132; 15'd10783: duty=135;
15'd10784: duty=136; 15'd10785: duty=143; 15'd10786: duty=135; 15'd10787: duty=128; 15'd10788: duty=132; 15'd10789: duty=129; 15'd10790: duty=125; 15'd10791: duty=128;
15'd10792: duty=121; 15'd10793: duty=113; 15'd10794: duty=113; 15'd10795: duty=114; 15'd10796: duty=120; 15'd10797: duty=114; 15'd10798: duty=107; 15'd10799: duty=112;
15'd10800: duty=113; 15'd10801: duty=111; 15'd10802: duty=113; 15'd10803: duty=107; 15'd10804: duty=110; 15'd10805: duty=116; 15'd10806: duty=118; 15'd10807: duty=116;
15'd10808: duty=115; 15'd10809: duty=119; 15'd10810: duty=114; 15'd10811: duty=112; 15'd10812: duty=118; 15'd10813: duty=107; 15'd10814: duty=99; 15'd10815: duty=108;
15'd10816: duty=107; 15'd10817: duty=113; 15'd10818: duty=115; 15'd10819: duty=118; 15'd10820: duty=116; 15'd10821: duty=117; 15'd10822: duty=118; 15'd10823: duty=124;
15'd10824: duty=131; 15'd10825: duty=129; 15'd10826: duty=127; 15'd10827: duty=125; 15'd10828: duty=134; 15'd10829: duty=135; 15'd10830: duty=127; 15'd10831: duty=132;
15'd10832: duty=141; 15'd10833: duty=145; 15'd10834: duty=148; 15'd10835: duty=149; 15'd10836: duty=145; 15'd10837: duty=146; 15'd10838: duty=147; 15'd10839: duty=143;
15'd10840: duty=144; 15'd10841: duty=142; 15'd10842: duty=145; 15'd10843: duty=142; 15'd10844: duty=151; 15'd10845: duty=159; 15'd10846: duty=157; 15'd10847: duty=160;
15'd10848: duty=156; 15'd10849: duty=161; 15'd10850: duty=159; 15'd10851: duty=156; 15'd10852: duty=151; 15'd10853: duty=153; 15'd10854: duty=149; 15'd10855: duty=142;
15'd10856: duty=148; 15'd10857: duty=153; 15'd10858: duty=145; 15'd10859: duty=139; 15'd10860: duty=143; 15'd10861: duty=147; 15'd10862: duty=145; 15'd10863: duty=139;
15'd10864: duty=132; 15'd10865: duty=126; 15'd10866: duty=122; 15'd10867: duty=117; 15'd10868: duty=113; 15'd10869: duty=125; 15'd10870: duty=128; 15'd10871: duty=116;
15'd10872: duty=116; 15'd10873: duty=110; 15'd10874: duty=116; 15'd10875: duty=123; 15'd10876: duty=111; 15'd10877: duty=98; 15'd10878: duty=102; 15'd10879: duty=105;
15'd10880: duty=105; 15'd10881: duty=96; 15'd10882: duty=96; 15'd10883: duty=98; 15'd10884: duty=104; 15'd10885: duty=104; 15'd10886: duty=106; 15'd10887: duty=110;
15'd10888: duty=107; 15'd10889: duty=116; 15'd10890: duty=110; 15'd10891: duty=122; 15'd10892: duty=124; 15'd10893: duty=121; 15'd10894: duty=122; 15'd10895: duty=116;
15'd10896: duty=118; 15'd10897: duty=126; 15'd10898: duty=125; 15'd10899: duty=122; 15'd10900: duty=134; 15'd10901: duty=137; 15'd10902: duty=131; 15'd10903: duty=133;
15'd10904: duty=133; 15'd10905: duty=139; 15'd10906: duty=136; 15'd10907: duty=140; 15'd10908: duty=138; 15'd10909: duty=139; 15'd10910: duty=141; 15'd10911: duty=139;
15'd10912: duty=145; 15'd10913: duty=149; 15'd10914: duty=159; 15'd10915: duty=153; 15'd10916: duty=157; 15'd10917: duty=153; 15'd10918: duty=151; 15'd10919: duty=154;
15'd10920: duty=159; 15'd10921: duty=160; 15'd10922: duty=159; 15'd10923: duty=153; 15'd10924: duty=151; 15'd10925: duty=155; 15'd10926: duty=157; 15'd10927: duty=153;
15'd10928: duty=142; 15'd10929: duty=145; 15'd10930: duty=137; 15'd10931: duty=132; 15'd10932: duty=143; 15'd10933: duty=140; 15'd10934: duty=135; 15'd10935: duty=143;
15'd10936: duty=134; 15'd10937: duty=134; 15'd10938: duty=139; 15'd10939: duty=142; 15'd10940: duty=144; 15'd10941: duty=139; 15'd10942: duty=134; 15'd10943: duty=127;
15'd10944: duty=125; 15'd10945: duty=119; 15'd10946: duty=113; 15'd10947: duty=112; 15'd10948: duty=108; 15'd10949: duty=101; 15'd10950: duty=111; 15'd10951: duty=115;
15'd10952: duty=115; 15'd10953: duty=113; 15'd10954: duty=103; 15'd10955: duty=106; 15'd10956: duty=99; 15'd10957: duty=95; 15'd10958: duty=96; 15'd10959: duty=97;
15'd10960: duty=102; 15'd10961: duty=101; 15'd10962: duty=102; 15'd10963: duty=104; 15'd10964: duty=109; 15'd10965: duty=113; 15'd10966: duty=112; 15'd10967: duty=114;
15'd10968: duty=118; 15'd10969: duty=110; 15'd10970: duty=105; 15'd10971: duty=116; 15'd10972: duty=113; 15'd10973: duty=125; 15'd10974: duty=128; 15'd10975: duty=128;
15'd10976: duty=136; 15'd10977: duty=131; 15'd10978: duty=134; 15'd10979: duty=131; 15'd10980: duty=137; 15'd10981: duty=136; 15'd10982: duty=136; 15'd10983: duty=139;
15'd10984: duty=142; 15'd10985: duty=144; 15'd10986: duty=151; 15'd10987: duty=157; 15'd10988: duty=162; 15'd10989: duty=160; 15'd10990: duty=152; 15'd10991: duty=154;
15'd10992: duty=163; 15'd10993: duty=168; 15'd10994: duty=164; 15'd10995: duty=161; 15'd10996: duty=160; 15'd10997: duty=162; 15'd10998: duty=158; 15'd10999: duty=151;
15'd11000: duty=151; 15'd11001: duty=146; 15'd11002: duty=145; 15'd11003: duty=150; 15'd11004: duty=142; 15'd11005: duty=146; 15'd11006: duty=141; 15'd11007: duty=140;
15'd11008: duty=129; 15'd11009: duty=129; 15'd11010: duty=139; 15'd11011: duty=140; 15'd11012: duty=145; 15'd11013: duty=149; 15'd11014: duty=141; 15'd11015: duty=134;
15'd11016: duty=135; 15'd11017: duty=132; 15'd11018: duty=128; 15'd11019: duty=129; 15'd11020: duty=123; 15'd11021: duty=123; 15'd11022: duty=112; 15'd11023: duty=100;
15'd11024: duty=103; 15'd11025: duty=96; 15'd11026: duty=105; 15'd11027: duty=96; 15'd11028: duty=105; 15'd11029: duty=108; 15'd11030: duty=107; 15'd11031: duty=116;
15'd11032: duty=106; 15'd11033: duty=116; 15'd11034: duty=115; 15'd11035: duty=103; 15'd11036: duty=100; 15'd11037: duty=92; 15'd11038: duty=98; 15'd11039: duty=103;
15'd11040: duty=106; 15'd11041: duty=107; 15'd11042: duty=112; 15'd11043: duty=121; 15'd11044: duty=118; 15'd11045: duty=114; 15'd11046: duty=118; 15'd11047: duty=129;
15'd11048: duty=123; 15'd11049: duty=132; 15'd11050: duty=131; 15'd11051: duty=132; 15'd11052: duty=130; 15'd11053: duty=124; 15'd11054: duty=123; 15'd11055: duty=113;
15'd11056: duty=127; 15'd11057: duty=146; 15'd11058: duty=147; 15'd11059: duty=142; 15'd11060: duty=147; 15'd11061: duty=146; 15'd11062: duty=151; 15'd11063: duty=151;
15'd11064: duty=150; 15'd11065: duty=154; 15'd11066: duty=164; 15'd11067: duty=173; 15'd11068: duty=168; 15'd11069: duty=165; 15'd11070: duty=156; 15'd11071: duty=157;
15'd11072: duty=156; 15'd11073: duty=156; 15'd11074: duty=156; 15'd11075: duty=151; 15'd11076: duty=147; 15'd11077: duty=148; 15'd11078: duty=154; 15'd11079: duty=146;
15'd11080: duty=150; 15'd11081: duty=153; 15'd11082: duty=157; 15'd11083: duty=154; 15'd11084: duty=148; 15'd11085: duty=145; 15'd11086: duty=134; 15'd11087: duty=139;
15'd11088: duty=136; 15'd11089: duty=121; 15'd11090: duty=133; 15'd11091: duty=134; 15'd11092: duty=122; 15'd11093: duty=123; 15'd11094: duty=122; 15'd11095: duty=130;
15'd11096: duty=125; 15'd11097: duty=115; 15'd11098: duty=110; 15'd11099: duty=124; 15'd11100: duty=127; 15'd11101: duty=116; 15'd11102: duty=111; 15'd11103: duty=102;
15'd11104: duty=94; 15'd11105: duty=100; 15'd11106: duty=103; 15'd11107: duty=104; 15'd11108: duty=102; 15'd11109: duty=104; 15'd11110: duty=118; 15'd11111: duty=118;
15'd11112: duty=112; 15'd11113: duty=103; 15'd11114: duty=105; 15'd11115: duty=100; 15'd11116: duty=107; 15'd11117: duty=101; 15'd11118: duty=104; 15'd11119: duty=104;
15'd11120: duty=108; 15'd11121: duty=119; 15'd11122: duty=124; 15'd11123: duty=128; 15'd11124: duty=121; 15'd11125: duty=121; 15'd11126: duty=121; 15'd11127: duty=127;
15'd11128: duty=121; 15'd11129: duty=118; 15'd11130: duty=121; 15'd11131: duty=127; 15'd11132: duty=130; 15'd11133: duty=132; 15'd11134: duty=135; 15'd11135: duty=132;
15'd11136: duty=128; 15'd11137: duty=138; 15'd11138: duty=145; 15'd11139: duty=160; 15'd11140: duty=162; 15'd11141: duty=166; 15'd11142: duty=165; 15'd11143: duty=166;
15'd11144: duty=170; 15'd11145: duty=156; 15'd11146: duty=161; 15'd11147: duty=157; 15'd11148: duty=145; 15'd11149: duty=149; 15'd11150: duty=159; 15'd11151: duty=165;
15'd11152: duty=170; 15'd11153: duty=173; 15'd11154: duty=162; 15'd11155: duty=148; 15'd11156: duty=159; 15'd11157: duty=163; 15'd11158: duty=155; 15'd11159: duty=157;
15'd11160: duty=154; 15'd11161: duty=158; 15'd11162: duty=153; 15'd11163: duty=146; 15'd11164: duty=150; 15'd11165: duty=134; 15'd11166: duty=141; 15'd11167: duty=137;
15'd11168: duty=128; 15'd11169: duty=133; 15'd11170: duty=134; 15'd11171: duty=121; 15'd11172: duty=120; 15'd11173: duty=111; 15'd11174: duty=99; 15'd11175: duty=116;
15'd11176: duty=96; 15'd11177: duty=104; 15'd11178: duty=107; 15'd11179: duty=101; 15'd11180: duty=99; 15'd11181: duty=92; 15'd11182: duty=101; 15'd11183: duty=93;
15'd11184: duty=101; 15'd11185: duty=102; 15'd11186: duty=96; 15'd11187: duty=104; 15'd11188: duty=107; 15'd11189: duty=101; 15'd11190: duty=85; 15'd11191: duty=102;
15'd11192: duty=102; 15'd11193: duty=92; 15'd11194: duty=98; 15'd11195: duty=99; 15'd11196: duty=105; 15'd11197: duty=96; 15'd11198: duty=105; 15'd11199: duty=115;
15'd11200: duty=126; 15'd11201: duty=128; 15'd11202: duty=122; 15'd11203: duty=130; 15'd11204: duty=134; 15'd11205: duty=137; 15'd11206: duty=134; 15'd11207: duty=131;
15'd11208: duty=126; 15'd11209: duty=125; 15'd11210: duty=135; 15'd11211: duty=137; 15'd11212: duty=139; 15'd11213: duty=140; 15'd11214: duty=135; 15'd11215: duty=146;
15'd11216: duty=153; 15'd11217: duty=151; 15'd11218: duty=145; 15'd11219: duty=152; 15'd11220: duty=164; 15'd11221: duty=165; 15'd11222: duty=175; 15'd11223: duty=174;
15'd11224: duty=164; 15'd11225: duty=174; 15'd11226: duty=173; 15'd11227: duty=172; 15'd11228: duty=168; 15'd11229: duty=157; 15'd11230: duty=165; 15'd11231: duty=160;
15'd11232: duty=159; 15'd11233: duty=159; 15'd11234: duty=153; 15'd11235: duty=155; 15'd11236: duty=151; 15'd11237: duty=142; 15'd11238: duty=147; 15'd11239: duty=137;
15'd11240: duty=134; 15'd11241: duty=146; 15'd11242: duty=137; 15'd11243: duty=131; 15'd11244: duty=139; 15'd11245: duty=140; 15'd11246: duty=126; 15'd11247: duty=118;
15'd11248: duty=118; 15'd11249: duty=119; 15'd11250: duty=124; 15'd11251: duty=123; 15'd11252: duty=114; 15'd11253: duty=107; 15'd11254: duty=111; 15'd11255: duty=110;
15'd11256: duty=111; 15'd11257: duty=106; 15'd11258: duty=105; 15'd11259: duty=106; 15'd11260: duty=104; 15'd11261: duty=112; 15'd11262: duty=102; 15'd11263: duty=102;
15'd11264: duty=97; 15'd11265: duty=93; 15'd11266: duty=105; 15'd11267: duty=104; 15'd11268: duty=110; 15'd11269: duty=108; 15'd11270: duty=109; 15'd11271: duty=129;
15'd11272: duty=117; 15'd11273: duty=119; 15'd11274: duty=117; 15'd11275: duty=112; 15'd11276: duty=129; 15'd11277: duty=121; 15'd11278: duty=113; 15'd11279: duty=108;
15'd11280: duty=112; 15'd11281: duty=117; 15'd11282: duty=117; 15'd11283: duty=112; 15'd11284: duty=113; 15'd11285: duty=112; 15'd11286: duty=129; 15'd11287: duty=127;
15'd11288: duty=129; 15'd11289: duty=131; 15'd11290: duty=131; 15'd11291: duty=138; 15'd11292: duty=143; 15'd11293: duty=141; 15'd11294: duty=143; 15'd11295: duty=156;
15'd11296: duty=154; 15'd11297: duty=154; 15'd11298: duty=151; 15'd11299: duty=156; 15'd11300: duty=159; 15'd11301: duty=165; 15'd11302: duty=159; 15'd11303: duty=155;
15'd11304: duty=156; 15'd11305: duty=159; 15'd11306: duty=159; 15'd11307: duty=152; 15'd11308: duty=147; 15'd11309: duty=155; 15'd11310: duty=155; 15'd11311: duty=162;
15'd11312: duty=158; 15'd11313: duty=160; 15'd11314: duty=158; 15'd11315: duty=158; 15'd11316: duty=159; 15'd11317: duty=158; 15'd11318: duty=156; 15'd11319: duty=144;
15'd11320: duty=135; 15'd11321: duty=131; 15'd11322: duty=138; 15'd11323: duty=139; 15'd11324: duty=138; 15'd11325: duty=132; 15'd11326: duty=141; 15'd11327: duty=132;
15'd11328: duty=126; 15'd11329: duty=128; 15'd11330: duty=113; 15'd11331: duty=105; 15'd11332: duty=115; 15'd11333: duty=110; 15'd11334: duty=123; 15'd11335: duty=107;
15'd11336: duty=112; 15'd11337: duty=110; 15'd11338: duty=107; 15'd11339: duty=102; 15'd11340: duty=96; 15'd11341: duty=115; 15'd11342: duty=98; 15'd11343: duty=95;
15'd11344: duty=103; 15'd11345: duty=99; 15'd11346: duty=95; 15'd11347: duty=96; 15'd11348: duty=96; 15'd11349: duty=108; 15'd11350: duty=106; 15'd11351: duty=96;
15'd11352: duty=83; 15'd11353: duty=96; 15'd11354: duty=106; 15'd11355: duty=107; 15'd11356: duty=106; 15'd11357: duty=119; 15'd11358: duty=124; 15'd11359: duty=124;
15'd11360: duty=131; 15'd11361: duty=132; 15'd11362: duty=127; 15'd11363: duty=135; 15'd11364: duty=144; 15'd11365: duty=135; 15'd11366: duty=135; 15'd11367: duty=132;
15'd11368: duty=123; 15'd11369: duty=123; 15'd11370: duty=136; 15'd11371: duty=140; 15'd11372: duty=148; 15'd11373: duty=146; 15'd11374: duty=147; 15'd11375: duty=148;
15'd11376: duty=146; 15'd11377: duty=146; 15'd11378: duty=152; 15'd11379: duty=154; 15'd11380: duty=156; 15'd11381: duty=154; 15'd11382: duty=155; 15'd11383: duty=161;
15'd11384: duty=167; 15'd11385: duty=168; 15'd11386: duty=173; 15'd11387: duty=168; 15'd11388: duty=165; 15'd11389: duty=168; 15'd11390: duty=169; 15'd11391: duty=160;
15'd11392: duty=158; 15'd11393: duty=162; 15'd11394: duty=156; 15'd11395: duty=162; 15'd11396: duty=162; 15'd11397: duty=153; 15'd11398: duty=145; 15'd11399: duty=151;
15'd11400: duty=146; 15'd11401: duty=143; 15'd11402: duty=134; 15'd11403: duty=128; 15'd11404: duty=130; 15'd11405: duty=125; 15'd11406: duty=121; 15'd11407: duty=118;
15'd11408: duty=113; 15'd11409: duty=110; 15'd11410: duty=101; 15'd11411: duty=109; 15'd11412: duty=118; 15'd11413: duty=112; 15'd11414: duty=121; 15'd11415: duty=112;
15'd11416: duty=106; 15'd11417: duty=119; 15'd11418: duty=113; 15'd11419: duty=105; 15'd11420: duty=98; 15'd11421: duty=94; 15'd11422: duty=96; 15'd11423: duty=102;
15'd11424: duty=109; 15'd11425: duty=109; 15'd11426: duty=107; 15'd11427: duty=97; 15'd11428: duty=108; 15'd11429: duty=117; 15'd11430: duty=116; 15'd11431: duty=113;
15'd11432: duty=104; 15'd11433: duty=113; 15'd11434: duty=117; 15'd11435: duty=107; 15'd11436: duty=103; 15'd11437: duty=97; 15'd11438: duty=109; 15'd11439: duty=112;
15'd11440: duty=114; 15'd11441: duty=127; 15'd11442: duty=128; 15'd11443: duty=119; 15'd11444: duty=121; 15'd11445: duty=113; 15'd11446: duty=124; 15'd11447: duty=138;
15'd11448: duty=124; 15'd11449: duty=111; 15'd11450: duty=118; 15'd11451: duty=131; 15'd11452: duty=138; 15'd11453: duty=149; 15'd11454: duty=147; 15'd11455: duty=146;
15'd11456: duty=145; 15'd11457: duty=152; 15'd11458: duty=153; 15'd11459: duty=156; 15'd11460: duty=159; 15'd11461: duty=162; 15'd11462: duty=160; 15'd11463: duty=171;
15'd11464: duty=165; 15'd11465: duty=164; 15'd11466: duty=173; 15'd11467: duty=167; 15'd11468: duty=163; 15'd11469: duty=164; 15'd11470: duty=160; 15'd11471: duty=161;
15'd11472: duty=157; 15'd11473: duty=154; 15'd11474: duty=149; 15'd11475: duty=158; 15'd11476: duty=163; 15'd11477: duty=162; 15'd11478: duty=163; 15'd11479: duty=159;
15'd11480: duty=151; 15'd11481: duty=144; 15'd11482: duty=149; 15'd11483: duty=141; 15'd11484: duty=137; 15'd11485: duty=127; 15'd11486: duty=127; 15'd11487: duty=118;
15'd11488: duty=127; 15'd11489: duty=126; 15'd11490: duty=128; 15'd11491: duty=117; 15'd11492: duty=116; 15'd11493: duty=124; 15'd11494: duty=119; 15'd11495: duty=115;
15'd11496: duty=116; 15'd11497: duty=106; 15'd11498: duty=102; 15'd11499: duty=115; 15'd11500: duty=111; 15'd11501: duty=105; 15'd11502: duty=94; 15'd11503: duty=92;
15'd11504: duty=87; 15'd11505: duty=104; 15'd11506: duty=100; 15'd11507: duty=86; 15'd11508: duty=88; 15'd11509: duty=98; 15'd11510: duty=103; 15'd11511: duty=103;
15'd11512: duty=111; 15'd11513: duty=109; 15'd11514: duty=103; 15'd11515: duty=115; 15'd11516: duty=114; 15'd11517: duty=120; 15'd11518: duty=119; 15'd11519: duty=115;
15'd11520: duty=114; 15'd11521: duty=120; 15'd11522: duty=124; 15'd11523: duty=116; 15'd11524: duty=121; 15'd11525: duty=121; 15'd11526: duty=122; 15'd11527: duty=128;
15'd11528: duty=131; 15'd11529: duty=134; 15'd11530: duty=136; 15'd11531: duty=131; 15'd11532: duty=132; 15'd11533: duty=139; 15'd11534: duty=148; 15'd11535: duty=145;
15'd11536: duty=153; 15'd11537: duty=154; 15'd11538: duty=149; 15'd11539: duty=153; 15'd11540: duty=154; 15'd11541: duty=157; 15'd11542: duty=162; 15'd11543: duty=165;
15'd11544: duty=163; 15'd11545: duty=162; 15'd11546: duty=168; 15'd11547: duty=163; 15'd11548: duty=159; 15'd11549: duty=162; 15'd11550: duty=168; 15'd11551: duty=177;
15'd11552: duty=173; 15'd11553: duty=179; 15'd11554: duty=168; 15'd11555: duty=154; 15'd11556: duty=151; 15'd11557: duty=147; 15'd11558: duty=146; 15'd11559: duty=136;
15'd11560: duty=140; 15'd11561: duty=139; 15'd11562: duty=136; 15'd11563: duty=137; 15'd11564: duty=130; 15'd11565: duty=136; 15'd11566: duty=136; 15'd11567: duty=127;
15'd11568: duty=121; 15'd11569: duty=127; 15'd11570: duty=122; 15'd11571: duty=107; 15'd11572: duty=108; 15'd11573: duty=99; 15'd11574: duty=96; 15'd11575: duty=109;
15'd11576: duty=108; 15'd11577: duty=113; 15'd11578: duty=113; 15'd11579: duty=113; 15'd11580: duty=110; 15'd11581: duty=104; 15'd11582: duty=105; 15'd11583: duty=106;
15'd11584: duty=105; 15'd11585: duty=101; 15'd11586: duty=102; 15'd11587: duty=106; 15'd11588: duty=112; 15'd11589: duty=109; 15'd11590: duty=107; 15'd11591: duty=112;
15'd11592: duty=118; 15'd11593: duty=102; 15'd11594: duty=93; 15'd11595: duty=92; 15'd11596: duty=98; 15'd11597: duty=110; 15'd11598: duty=125; 15'd11599: duty=123;
15'd11600: duty=119; 15'd11601: duty=119; 15'd11602: duty=127; 15'd11603: duty=127; 15'd11604: duty=121; 15'd11605: duty=123; 15'd11606: duty=124; 15'd11607: duty=127;
15'd11608: duty=127; 15'd11609: duty=131; 15'd11610: duty=126; 15'd11611: duty=128; 15'd11612: duty=138; 15'd11613: duty=141; 15'd11614: duty=138; 15'd11615: duty=145;
15'd11616: duty=147; 15'd11617: duty=149; 15'd11618: duty=153; 15'd11619: duty=155; 15'd11620: duty=144; 15'd11621: duty=152; 15'd11622: duty=159; 15'd11623: duty=158;
15'd11624: duty=161; 15'd11625: duty=161; 15'd11626: duty=160; 15'd11627: duty=161; 15'd11628: duty=156; 15'd11629: duty=158; 15'd11630: duty=161; 15'd11631: duty=165;
15'd11632: duty=170; 15'd11633: duty=172; 15'd11634: duty=174; 15'd11635: duty=169; 15'd11636: duty=164; 15'd11637: duty=159; 15'd11638: duty=152; 15'd11639: duty=144;
15'd11640: duty=146; 15'd11641: duty=141; 15'd11642: duty=142; 15'd11643: duty=141; 15'd11644: duty=138; 15'd11645: duty=133; 15'd11646: duty=127; 15'd11647: duty=126;
15'd11648: duty=132; 15'd11649: duty=131; 15'd11650: duty=128; 15'd11651: duty=118; 15'd11652: duty=122; 15'd11653: duty=128; 15'd11654: duty=127; 15'd11655: duty=120;
15'd11656: duty=106; 15'd11657: duty=102; 15'd11658: duty=109; 15'd11659: duty=109; 15'd11660: duty=106; 15'd11661: duty=99; 15'd11662: duty=99; 15'd11663: duty=116;
15'd11664: duty=119; 15'd11665: duty=113; 15'd11666: duty=101; 15'd11667: duty=104; 15'd11668: duty=104; 15'd11669: duty=109; 15'd11670: duty=104; 15'd11671: duty=103;
15'd11672: duty=99; 15'd11673: duty=92; 15'd11674: duty=108; 15'd11675: duty=114; 15'd11676: duty=108; 15'd11677: duty=106; 15'd11678: duty=110; 15'd11679: duty=113;
15'd11680: duty=114; 15'd11681: duty=117; 15'd11682: duty=113; 15'd11683: duty=114; 15'd11684: duty=112; 15'd11685: duty=111; 15'd11686: duty=117; 15'd11687: duty=122;
15'd11688: duty=123; 15'd11689: duty=126; 15'd11690: duty=122; 15'd11691: duty=122; 15'd11692: duty=132; 15'd11693: duty=135; 15'd11694: duty=136; 15'd11695: duty=126;
15'd11696: duty=129; 15'd11697: duty=143; 15'd11698: duty=144; 15'd11699: duty=143; 15'd11700: duty=138; 15'd11701: duty=138; 15'd11702: duty=150; 15'd11703: duty=164;
15'd11704: duty=160; 15'd11705: duty=161; 15'd11706: duty=167; 15'd11707: duty=159; 15'd11708: duty=169; 15'd11709: duty=166; 15'd11710: duty=169; 15'd11711: duty=178;
15'd11712: duty=169; 15'd11713: duty=162; 15'd11714: duty=162; 15'd11715: duty=165; 15'd11716: duty=163; 15'd11717: duty=170; 15'd11718: duty=163; 15'd11719: duty=159;
15'd11720: duty=157; 15'd11721: duty=159; 15'd11722: duty=157; 15'd11723: duty=153; 15'd11724: duty=156; 15'd11725: duty=145; 15'd11726: duty=141; 15'd11727: duty=136;
15'd11728: duty=145; 15'd11729: duty=139; 15'd11730: duty=127; 15'd11731: duty=124; 15'd11732: duty=119; 15'd11733: duty=125; 15'd11734: duty=126; 15'd11735: duty=114;
15'd11736: duty=110; 15'd11737: duty=107; 15'd11738: duty=104; 15'd11739: duty=114; 15'd11740: duty=108; 15'd11741: duty=107; 15'd11742: duty=109; 15'd11743: duty=105;
15'd11744: duty=104; 15'd11745: duty=107; 15'd11746: duty=101; 15'd11747: duty=99; 15'd11748: duty=106; 15'd11749: duty=108; 15'd11750: duty=103; 15'd11751: duty=102;
15'd11752: duty=92; 15'd11753: duty=91; 15'd11754: duty=101; 15'd11755: duty=110; 15'd11756: duty=107; 15'd11757: duty=110; 15'd11758: duty=113; 15'd11759: duty=111;
15'd11760: duty=106; 15'd11761: duty=107; 15'd11762: duty=112; 15'd11763: duty=122; 15'd11764: duty=123; 15'd11765: duty=122; 15'd11766: duty=120; 15'd11767: duty=114;
15'd11768: duty=113; 15'd11769: duty=117; 15'd11770: duty=138; 15'd11771: duty=143; 15'd11772: duty=139; 15'd11773: duty=125; 15'd11774: duty=127; 15'd11775: duty=124;
15'd11776: duty=123; 15'd11777: duty=127; 15'd11778: duty=127; 15'd11779: duty=132; 15'd11780: duty=138; 15'd11781: duty=140; 15'd11782: duty=153; 15'd11783: duty=151;
15'd11784: duty=152; 15'd11785: duty=149; 15'd11786: duty=151; 15'd11787: duty=160; 15'd11788: duty=159; 15'd11789: duty=160; 15'd11790: duty=154; 15'd11791: duty=152;
15'd11792: duty=150; 15'd11793: duty=151; 15'd11794: duty=155; 15'd11795: duty=156; 15'd11796: duty=165; 15'd11797: duty=163; 15'd11798: duty=167; 15'd11799: duty=165;
15'd11800: duty=162; 15'd11801: duty=174; 15'd11802: duty=163; 15'd11803: duty=162; 15'd11804: duty=160; 15'd11805: duty=156; 15'd11806: duty=147; 15'd11807: duty=157;
15'd11808: duty=151; 15'd11809: duty=143; 15'd11810: duty=145; 15'd11811: duty=142; 15'd11812: duty=137; 15'd11813: duty=133; 15'd11814: duty=128; 15'd11815: duty=139;
15'd11816: duty=136; 15'd11817: duty=131; 15'd11818: duty=124; 15'd11819: duty=104; 15'd11820: duty=115; 15'd11821: duty=118; 15'd11822: duty=121; 15'd11823: duty=124;
15'd11824: duty=110; 15'd11825: duty=112; 15'd11826: duty=108; 15'd11827: duty=96; 15'd11828: duty=108; 15'd11829: duty=104; 15'd11830: duty=102; 15'd11831: duty=101;
15'd11832: duty=98; 15'd11833: duty=95; 15'd11834: duty=96; 15'd11835: duty=102; 15'd11836: duty=104; 15'd11837: duty=109; 15'd11838: duty=108; 15'd11839: duty=103;
15'd11840: duty=99; 15'd11841: duty=92; 15'd11842: duty=101; 15'd11843: duty=108; 15'd11844: duty=108; 15'd11845: duty=105; 15'd11846: duty=110; 15'd11847: duty=125;
15'd11848: duty=127; 15'd11849: duty=127; 15'd11850: duty=127; 15'd11851: duty=128; 15'd11852: duty=129; 15'd11853: duty=125; 15'd11854: duty=129; 15'd11855: duty=127;
15'd11856: duty=119; 15'd11857: duty=115; 15'd11858: duty=128; 15'd11859: duty=131; 15'd11860: duty=137; 15'd11861: duty=147; 15'd11862: duty=134; 15'd11863: duty=140;
15'd11864: duty=150; 15'd11865: duty=147; 15'd11866: duty=150; 15'd11867: duty=150; 15'd11868: duty=150; 15'd11869: duty=157; 15'd11870: duty=157; 15'd11871: duty=151;
15'd11872: duty=150; 15'd11873: duty=151; 15'd11874: duty=150; 15'd11875: duty=157; 15'd11876: duty=162; 15'd11877: duty=156; 15'd11878: duty=148; 15'd11879: duty=154;
15'd11880: duty=154; 15'd11881: duty=153; 15'd11882: duty=154; 15'd11883: duty=156; 15'd11884: duty=158; 15'd11885: duty=171; 15'd11886: duty=168; 15'd11887: duty=163;
15'd11888: duty=168; 15'd11889: duty=162; 15'd11890: duty=157; 15'd11891: duty=154; 15'd11892: duty=151; 15'd11893: duty=146; 15'd11894: duty=148; 15'd11895: duty=137;
15'd11896: duty=137; 15'd11897: duty=133; 15'd11898: duty=131; 15'd11899: duty=133; 15'd11900: duty=124; 15'd11901: duty=119; 15'd11902: duty=119; 15'd11903: duty=112;
15'd11904: duty=114; 15'd11905: duty=116; 15'd11906: duty=118; 15'd11907: duty=119; 15'd11908: duty=110; 15'd11909: duty=106; 15'd11910: duty=102; 15'd11911: duty=98;
15'd11912: duty=96; 15'd11913: duty=95; 15'd11914: duty=101; 15'd11915: duty=101; 15'd11916: duty=98; 15'd11917: duty=92; 15'd11918: duty=96; 15'd11919: duty=102;
15'd11920: duty=96; 15'd11921: duty=110; 15'd11922: duty=104; 15'd11923: duty=112; 15'd11924: duty=124; 15'd11925: duty=119; 15'd11926: duty=111; 15'd11927: duty=105;
15'd11928: duty=116; 15'd11929: duty=119; 15'd11930: duty=121; 15'd11931: duty=113; 15'd11932: duty=118; 15'd11933: duty=121; 15'd11934: duty=124; 15'd11935: duty=132;
15'd11936: duty=125; 15'd11937: duty=121; 15'd11938: duty=122; 15'd11939: duty=124; 15'd11940: duty=121; 15'd11941: duty=114; 15'd11942: duty=119; 15'd11943: duty=127;
15'd11944: duty=130; 15'd11945: duty=133; 15'd11946: duty=126; 15'd11947: duty=137; 15'd11948: duty=145; 15'd11949: duty=151; 15'd11950: duty=159; 15'd11951: duty=153;
15'd11952: duty=157; 15'd11953: duty=155; 15'd11954: duty=156; 15'd11955: duty=166; 15'd11956: duty=163; 15'd11957: duty=152; 15'd11958: duty=154; 15'd11959: duty=154;
15'd11960: duty=153; 15'd11961: duty=162; 15'd11962: duty=159; 15'd11963: duty=159; 15'd11964: duty=154; 15'd11965: duty=149; 15'd11966: duty=156; 15'd11967: duty=156;
15'd11968: duty=154; 15'd11969: duty=150; 15'd11970: duty=157; 15'd11971: duty=157; 15'd11972: duty=162; 15'd11973: duty=154; 15'd11974: duty=156; 15'd11975: duty=157;
15'd11976: duty=147; 15'd11977: duty=145; 15'd11978: duty=145; 15'd11979: duty=142; 15'd11980: duty=134; 15'd11981: duty=136; 15'd11982: duty=129; 15'd11983: duty=125;
15'd11984: duty=128; 15'd11985: duty=126; 15'd11986: duty=114; 15'd11987: duty=113; 15'd11988: duty=116; 15'd11989: duty=115; 15'd11990: duty=113; 15'd11991: duty=113;
15'd11992: duty=108; 15'd11993: duty=113; 15'd11994: duty=116; 15'd11995: duty=109; 15'd11996: duty=102; 15'd11997: duty=99; 15'd11998: duty=107; 15'd11999: duty=107;
15'd12000: duty=107; 15'd12001: duty=112; 15'd12002: duty=111; 15'd12003: duty=104; 15'd12004: duty=104; 15'd12005: duty=107; 15'd12006: duty=107; 15'd12007: duty=108;
15'd12008: duty=107; 15'd12009: duty=112; 15'd12010: duty=116; 15'd12011: duty=115; 15'd12012: duty=103; 15'd12013: duty=101; 15'd12014: duty=113; 15'd12015: duty=107;
15'd12016: duty=111; 15'd12017: duty=120; 15'd12018: duty=121; 15'd12019: duty=120; 15'd12020: duty=123; 15'd12021: duty=126; 15'd12022: duty=119; 15'd12023: duty=123;
15'd12024: duty=131; 15'd12025: duty=133; 15'd12026: duty=128; 15'd12027: duty=123; 15'd12028: duty=135; 15'd12029: duty=138; 15'd12030: duty=127; 15'd12031: duty=130;
15'd12032: duty=140; 15'd12033: duty=137; 15'd12034: duty=142; 15'd12035: duty=159; 15'd12036: duty=143; 15'd12037: duty=138; 15'd12038: duty=145; 15'd12039: duty=148;
15'd12040: duty=154; 15'd12041: duty=150; 15'd12042: duty=156; 15'd12043: duty=153; 15'd12044: duty=153; 15'd12045: duty=158; 15'd12046: duty=160; 15'd12047: duty=160;
15'd12048: duty=163; 15'd12049: duty=163; 15'd12050: duty=165; 15'd12051: duty=159; 15'd12052: duty=160; 15'd12053: duty=165; 15'd12054: duty=160; 15'd12055: duty=162;
15'd12056: duty=166; 15'd12057: duty=162; 15'd12058: duty=159; 15'd12059: duty=154; 15'd12060: duty=154; 15'd12061: duty=153; 15'd12062: duty=146; 15'd12063: duty=144;
15'd12064: duty=142; 15'd12065: duty=139; 15'd12066: duty=129; 15'd12067: duty=125; 15'd12068: duty=124; 15'd12069: duty=124; 15'd12070: duty=124; 15'd12071: duty=129;
15'd12072: duty=124; 15'd12073: duty=113; 15'd12074: duty=116; 15'd12075: duty=116; 15'd12076: duty=108; 15'd12077: duty=107; 15'd12078: duty=105; 15'd12079: duty=102;
15'd12080: duty=102; 15'd12081: duty=101; 15'd12082: duty=95; 15'd12083: duty=101; 15'd12084: duty=102; 15'd12085: duty=99; 15'd12086: duty=107; 15'd12087: duty=101;
15'd12088: duty=96; 15'd12089: duty=101; 15'd12090: duty=98; 15'd12091: duty=98; 15'd12092: duty=107; 15'd12093: duty=110; 15'd12094: duty=113; 15'd12095: duty=113;
15'd12096: duty=107; 15'd12097: duty=101; 15'd12098: duty=111; 15'd12099: duty=113; 15'd12100: duty=119; 15'd12101: duty=128; 15'd12102: duty=131; 15'd12103: duty=130;
15'd12104: duty=118; 15'd12105: duty=110; 15'd12106: duty=116; 15'd12107: duty=124; 15'd12108: duty=124; 15'd12109: duty=131; 15'd12110: duty=127; 15'd12111: duty=131;
15'd12112: duty=134; 15'd12113: duty=130; 15'd12114: duty=131; 15'd12115: duty=124; 15'd12116: duty=139; 15'd12117: duty=133; 15'd12118: duty=133; 15'd12119: duty=134;
15'd12120: duty=134; 15'd12121: duty=144; 15'd12122: duty=148; 15'd12123: duty=147; 15'd12124: duty=148; 15'd12125: duty=151; 15'd12126: duty=151; 15'd12127: duty=168;
15'd12128: duty=157; 15'd12129: duty=153; 15'd12130: duty=163; 15'd12131: duty=164; 15'd12132: duty=163; 15'd12133: duty=160; 15'd12134: duty=156; 15'd12135: duty=157;
15'd12136: duty=156; 15'd12137: duty=161; 15'd12138: duty=157; 15'd12139: duty=157; 15'd12140: duty=159; 15'd12141: duty=162; 15'd12142: duty=161; 15'd12143: duty=162;
15'd12144: duty=157; 15'd12145: duty=153; 15'd12146: duty=155; 15'd12147: duty=147; 15'd12148: duty=144; 15'd12149: duty=143; 15'd12150: duty=145; 15'd12151: duty=146;
15'd12152: duty=147; 15'd12153: duty=146; 15'd12154: duty=137; 15'd12155: duty=134; 15'd12156: duty=126; 15'd12157: duty=121; 15'd12158: duty=119; 15'd12159: duty=116;
15'd12160: duty=115; 15'd12161: duty=110; 15'd12162: duty=107; 15'd12163: duty=107; 15'd12164: duty=111; 15'd12165: duty=108; 15'd12166: duty=113; 15'd12167: duty=107;
15'd12168: duty=101; 15'd12169: duty=99; 15'd12170: duty=104; 15'd12171: duty=99; 15'd12172: duty=105; 15'd12173: duty=99; 15'd12174: duty=99; 15'd12175: duty=99;
15'd12176: duty=98; 15'd12177: duty=110; 15'd12178: duty=110; 15'd12179: duty=108; 15'd12180: duty=103; 15'd12181: duty=108; 15'd12182: duty=107; 15'd12183: duty=108;
15'd12184: duty=109; 15'd12185: duty=108; 15'd12186: duty=106; 15'd12187: duty=107; 15'd12188: duty=106; 15'd12189: duty=116; 15'd12190: duty=124; 15'd12191: duty=127;
15'd12192: duty=131; 15'd12193: duty=128; 15'd12194: duty=123; 15'd12195: duty=127; 15'd12196: duty=124; 15'd12197: duty=128; 15'd12198: duty=126; 15'd12199: duty=129;
15'd12200: duty=124; 15'd12201: duty=124; 15'd12202: duty=129; 15'd12203: duty=131; 15'd12204: duty=134; 15'd12205: duty=132; 15'd12206: duty=133; 15'd12207: duty=143;
15'd12208: duty=147; 15'd12209: duty=143; 15'd12210: duty=151; 15'd12211: duty=149; 15'd12212: duty=151; 15'd12213: duty=156; 15'd12214: duty=154; 15'd12215: duty=149;
15'd12216: duty=153; 15'd12217: duty=153; 15'd12218: duty=161; 15'd12219: duty=163; 15'd12220: duty=166; 15'd12221: duty=166; 15'd12222: duty=160; 15'd12223: duty=154;
15'd12224: duty=168; 15'd12225: duty=166; 15'd12226: duty=168; 15'd12227: duty=163; 15'd12228: duty=149; 15'd12229: duty=147; 15'd12230: duty=149; 15'd12231: duty=156;
15'd12232: duty=157; 15'd12233: duty=162; 15'd12234: duty=157; 15'd12235: duty=162; 15'd12236: duty=154; 15'd12237: duty=154; 15'd12238: duty=146; 15'd12239: duty=134;
15'd12240: duty=132; 15'd12241: duty=139; 15'd12242: duty=142; 15'd12243: duty=141; 15'd12244: duty=136; 15'd12245: duty=126; 15'd12246: duty=119; 15'd12247: duty=118;
15'd12248: duty=121; 15'd12249: duty=118; 15'd12250: duty=114; 15'd12251: duty=104; 15'd12252: duty=108; 15'd12253: duty=114; 15'd12254: duty=108; 15'd12255: duty=106;
15'd12256: duty=103; 15'd12257: duty=99; 15'd12258: duty=102; 15'd12259: duty=105; 15'd12260: duty=97; 15'd12261: duty=93; 15'd12262: duty=94; 15'd12263: duty=98;
15'd12264: duty=97; 15'd12265: duty=95; 15'd12266: duty=96; 15'd12267: duty=96; 15'd12268: duty=99; 15'd12269: duty=107; 15'd12270: duty=107; 15'd12271: duty=105;
15'd12272: duty=109; 15'd12273: duty=101; 15'd12274: duty=107; 15'd12275: duty=113; 15'd12276: duty=112; 15'd12277: duty=106; 15'd12278: duty=107; 15'd12279: duty=115;
15'd12280: duty=120; 15'd12281: duty=125; 15'd12282: duty=134; 15'd12283: duty=132; 15'd12284: duty=131; 15'd12285: duty=134; 15'd12286: duty=134; 15'd12287: duty=136;
15'd12288: duty=124; 15'd12289: duty=126; 15'd12290: duty=134; 15'd12291: duty=134; 15'd12292: duty=140; 15'd12293: duty=137; 15'd12294: duty=133; 15'd12295: duty=139;
15'd12296: duty=145; 15'd12297: duty=150; 15'd12298: duty=148; 15'd12299: duty=157; 15'd12300: duty=151; 15'd12301: duty=154; 15'd12302: duty=156; 15'd12303: duty=150;
15'd12304: duty=152; 15'd12305: duty=154; 15'd12306: duty=160; 15'd12307: duty=160; 15'd12308: duty=163; 15'd12309: duty=160; 15'd12310: duty=162; 15'd12311: duty=165;
15'd12312: duty=161; 15'd12313: duty=162; 15'd12314: duty=165; 15'd12315: duty=165; 15'd12316: duty=173; 15'd12317: duty=168; 15'd12318: duty=161; 15'd12319: duty=163;
15'd12320: duty=164; 15'd12321: duty=156; 15'd12322: duty=150; 15'd12323: duty=143; 15'd12324: duty=146; 15'd12325: duty=148; 15'd12326: duty=144; 15'd12327: duty=142;
15'd12328: duty=131; 15'd12329: duty=131; 15'd12330: duty=133; 15'd12331: duty=134; 15'd12332: duty=133; 15'd12333: duty=131; 15'd12334: duty=126; 15'd12335: duty=127;
15'd12336: duty=112; 15'd12337: duty=105; 15'd12338: duty=109; 15'd12339: duty=106; 15'd12340: duty=105; 15'd12341: duty=106; 15'd12342: duty=96; 15'd12343: duty=97;
15'd12344: duty=101; 15'd12345: duty=97; 15'd12346: duty=105; 15'd12347: duty=105; 15'd12348: duty=105; 15'd12349: duty=105; 15'd12350: duty=104; 15'd12351: duty=102;
15'd12352: duty=104; 15'd12353: duty=101; 15'd12354: duty=104; 15'd12355: duty=105; 15'd12356: duty=103; 15'd12357: duty=107; 15'd12358: duty=107; 15'd12359: duty=103;
15'd12360: duty=98; 15'd12361: duty=103; 15'd12362: duty=104; 15'd12363: duty=110; 15'd12364: duty=106; 15'd12365: duty=104; 15'd12366: duty=113; 15'd12367: duty=113;
15'd12368: duty=121; 15'd12369: duty=124; 15'd12370: duty=118; 15'd12371: duty=124; 15'd12372: duty=127; 15'd12373: duty=130; 15'd12374: duty=139; 15'd12375: duty=136;
15'd12376: duty=128; 15'd12377: duty=128; 15'd12378: duty=131; 15'd12379: duty=132; 15'd12380: duty=133; 15'd12381: duty=134; 15'd12382: duty=136; 15'd12383: duty=139;
15'd12384: duty=149; 15'd12385: duty=149; 15'd12386: duty=150; 15'd12387: duty=143; 15'd12388: duty=137; 15'd12389: duty=146; 15'd12390: duty=147; 15'd12391: duty=156;
15'd12392: duty=155; 15'd12393: duty=149; 15'd12394: duty=154; 15'd12395: duty=162; 15'd12396: duty=165; 15'd12397: duty=160; 15'd12398: duty=156; 15'd12399: duty=165;
15'd12400: duty=164; 15'd12401: duty=162; 15'd12402: duty=167; 15'd12403: duty=164; 15'd12404: duty=153; 15'd12405: duty=151; 15'd12406: duty=160; 15'd12407: duty=159;
15'd12408: duty=157; 15'd12409: duty=162; 15'd12410: duty=159; 15'd12411: duty=158; 15'd12412: duty=154; 15'd12413: duty=148; 15'd12414: duty=150; 15'd12415: duty=151;
15'd12416: duty=154; 15'd12417: duty=148; 15'd12418: duty=146; 15'd12419: duty=145; 15'd12420: duty=145; 15'd12421: duty=142; 15'd12422: duty=137; 15'd12423: duty=130;
15'd12424: duty=133; 15'd12425: duty=131; 15'd12426: duty=121; 15'd12427: duty=121; 15'd12428: duty=110; 15'd12429: duty=105; 15'd12430: duty=110; 15'd12431: duty=104;
15'd12432: duty=97; 15'd12433: duty=99; 15'd12434: duty=94; 15'd12435: duty=92; 15'd12436: duty=91; 15'd12437: duty=94; 15'd12438: duty=93; 15'd12439: duty=91;
15'd12440: duty=88; 15'd12441: duty=85; 15'd12442: duty=91; 15'd12443: duty=92; 15'd12444: duty=98; 15'd12445: duty=95; 15'd12446: duty=99; 15'd12447: duty=106;
15'd12448: duty=110; 15'd12449: duty=111; 15'd12450: duty=107; 15'd12451: duty=110; 15'd12452: duty=111; 15'd12453: duty=107; 15'd12454: duty=110; 15'd12455: duty=118;
15'd12456: duty=110; 15'd12457: duty=117; 15'd12458: duty=127; 15'd12459: duty=125; 15'd12460: duty=131; 15'd12461: duty=131; 15'd12462: duty=121; 15'd12463: duty=122;
15'd12464: duty=130; 15'd12465: duty=128; 15'd12466: duty=130; 15'd12467: duty=132; 15'd12468: duty=130; 15'd12469: duty=139; 15'd12470: duty=136; 15'd12471: duty=140;
15'd12472: duty=136; 15'd12473: duty=134; 15'd12474: duty=147; 15'd12475: duty=145; 15'd12476: duty=144; 15'd12477: duty=143; 15'd12478: duty=150; 15'd12479: duty=154;
15'd12480: duty=154; 15'd12481: duty=154; 15'd12482: duty=158; 15'd12483: duty=154; 15'd12484: duty=148; 15'd12485: duty=149; 15'd12486: duty=157; 15'd12487: duty=165;
15'd12488: duty=163; 15'd12489: duty=162; 15'd12490: duty=158; 15'd12491: duty=153; 15'd12492: duty=157; 15'd12493: duty=159; 15'd12494: duty=159; 15'd12495: duty=164;
15'd12496: duty=165; 15'd12497: duty=164; 15'd12498: duty=166; 15'd12499: duty=162; 15'd12500: duty=152; 15'd12501: duty=153; 15'd12502: duty=154; 15'd12503: duty=148;
15'd12504: duty=153; 15'd12505: duty=161; 15'd12506: duty=154; 15'd12507: duty=150; 15'd12508: duty=140; 15'd12509: duty=133; 15'd12510: duty=139; 15'd12511: duty=133;
15'd12512: duty=127; 15'd12513: duty=122; 15'd12514: duty=123; 15'd12515: duty=121; 15'd12516: duty=115; 15'd12517: duty=115; 15'd12518: duty=107; 15'd12519: duty=108;
15'd12520: duty=107; 15'd12521: duty=111; 15'd12522: duty=109; 15'd12523: duty=101; 15'd12524: duty=96; 15'd12525: duty=93; 15'd12526: duty=93; 15'd12527: duty=97;
15'd12528: duty=101; 15'd12529: duty=98; 15'd12530: duty=93; 15'd12531: duty=93; 15'd12532: duty=95; 15'd12533: duty=99; 15'd12534: duty=102; 15'd12535: duty=105;
15'd12536: duty=105; 15'd12537: duty=97; 15'd12538: duty=101; 15'd12539: duty=104; 15'd12540: duty=107; 15'd12541: duty=110; 15'd12542: duty=113; 15'd12543: duty=116;
15'd12544: duty=118; 15'd12545: duty=124; 15'd12546: duty=126; 15'd12547: duty=122; 15'd12548: duty=123; 15'd12549: duty=127; 15'd12550: duty=131; 15'd12551: duty=122;
15'd12552: duty=115; 15'd12553: duty=117; 15'd12554: duty=126; 15'd12555: duty=138; 15'd12556: duty=133; 15'd12557: duty=137; 15'd12558: duty=130; 15'd12559: duty=134;
15'd12560: duty=148; 15'd12561: duty=139; 15'd12562: duty=136; 15'd12563: duty=142; 15'd12564: duty=142; 15'd12565: duty=141; 15'd12566: duty=144; 15'd12567: duty=157;
15'd12568: duty=145; 15'd12569: duty=142; 15'd12570: duty=155; 15'd12571: duty=143; 15'd12572: duty=136; 15'd12573: duty=151; 15'd12574: duty=153; 15'd12575: duty=150;
15'd12576: duty=153; 15'd12577: duty=153; 15'd12578: duty=153; 15'd12579: duty=154; 15'd12580: duty=167; 15'd12581: duty=162; 15'd12582: duty=166; 15'd12583: duty=160;
15'd12584: duty=156; 15'd12585: duty=162; 15'd12586: duty=159; 15'd12587: duty=157; 15'd12588: duty=159; 15'd12589: duty=160; 15'd12590: duty=160; 15'd12591: duty=160;
15'd12592: duty=159; 15'd12593: duty=161; 15'd12594: duty=158; 15'd12595: duty=160; 15'd12596: duty=157; 15'd12597: duty=150; 15'd12598: duty=153; 15'd12599: duty=149;
15'd12600: duty=142; 15'd12601: duty=142; 15'd12602: duty=139; 15'd12603: duty=127; 15'd12604: duty=121; 15'd12605: duty=116; 15'd12606: duty=112; 15'd12607: duty=113;
15'd12608: duty=110; 15'd12609: duty=107; 15'd12610: duty=102; 15'd12611: duty=96; 15'd12612: duty=96; 15'd12613: duty=95; 15'd12614: duty=87; 15'd12615: duty=96;
15'd12616: duty=93; 15'd12617: duty=92; 15'd12618: duty=92; 15'd12619: duty=82; 15'd12620: duty=80; 15'd12621: duty=87; 15'd12622: duty=87; 15'd12623: duty=96;
15'd12624: duty=102; 15'd12625: duty=103; 15'd12626: duty=106; 15'd12627: duty=108; 15'd12628: duty=105; 15'd12629: duty=111; 15'd12630: duty=110; 15'd12631: duty=102;
15'd12632: duty=109; 15'd12633: duty=114; 15'd12634: duty=113; 15'd12635: duty=113; 15'd12636: duty=115; 15'd12637: duty=118; 15'd12638: duty=130; 15'd12639: duty=132;
15'd12640: duty=137; 15'd12641: duty=131; 15'd12642: duty=124; 15'd12643: duty=133; 15'd12644: duty=139; 15'd12645: duty=131; 15'd12646: duty=130; 15'd12647: duty=128;
15'd12648: duty=139; 15'd12649: duty=141; 15'd12650: duty=140; 15'd12651: duty=136; 15'd12652: duty=133; 15'd12653: duty=145; 15'd12654: duty=147; 15'd12655: duty=151;
15'd12656: duty=148; 15'd12657: duty=148; 15'd12658: duty=145; 15'd12659: duty=148; 15'd12660: duty=160; 15'd12661: duty=165; 15'd12662: duty=157; 15'd12663: duty=156;
15'd12664: duty=165; 15'd12665: duty=165; 15'd12666: duty=167; 15'd12667: duty=167; 15'd12668: duty=161; 15'd12669: duty=170; 15'd12670: duty=167; 15'd12671: duty=163;
15'd12672: duty=156; 15'd12673: duty=151; 15'd12674: duty=151; 15'd12675: duty=151; 15'd12676: duty=157; 15'd12677: duty=156; 15'd12678: duty=157; 15'd12679: duty=151;
15'd12680: duty=151; 15'd12681: duty=154; 15'd12682: duty=151; 15'd12683: duty=153; 15'd12684: duty=145; 15'd12685: duty=145; 15'd12686: duty=148; 15'd12687: duty=149;
15'd12688: duty=147; 15'd12689: duty=137; 15'd12690: duty=133; 15'd12691: duty=127; 15'd12692: duty=119; 15'd12693: duty=124; 15'd12694: duty=113; 15'd12695: duty=106;
15'd12696: duty=107; 15'd12697: duty=104; 15'd12698: duty=104; 15'd12699: duty=98; 15'd12700: duty=98; 15'd12701: duty=92; 15'd12702: duty=95; 15'd12703: duty=95;
15'd12704: duty=104; 15'd12705: duty=101; 15'd12706: duty=98; 15'd12707: duty=98; 15'd12708: duty=99; 15'd12709: duty=105; 15'd12710: duty=99; 15'd12711: duty=99;
15'd12712: duty=96; 15'd12713: duty=106; 15'd12714: duty=107; 15'd12715: duty=107; 15'd12716: duty=107; 15'd12717: duty=103; 15'd12718: duty=110; 15'd12719: duty=96;
15'd12720: duty=99; 15'd12721: duty=109; 15'd12722: duty=105; 15'd12723: duty=107; 15'd12724: duty=116; 15'd12725: duty=118; 15'd12726: duty=119; 15'd12727: duty=121;
15'd12728: duty=120; 15'd12729: duty=118; 15'd12730: duty=119; 15'd12731: duty=133; 15'd12732: duty=125; 15'd12733: duty=124; 15'd12734: duty=136; 15'd12735: duty=130;
15'd12736: duty=128; 15'd12737: duty=137; 15'd12738: duty=139; 15'd12739: duty=148; 15'd12740: duty=142; 15'd12741: duty=139; 15'd12742: duty=148; 15'd12743: duty=142;
15'd12744: duty=153; 15'd12745: duty=163; 15'd12746: duty=159; 15'd12747: duty=156; 15'd12748: duty=149; 15'd12749: duty=159; 15'd12750: duty=162; 15'd12751: duty=151;
15'd12752: duty=160; 15'd12753: duty=161; 15'd12754: duty=148; 15'd12755: duty=150; 15'd12756: duty=158; 15'd12757: duty=162; 15'd12758: duty=164; 15'd12759: duty=159;
15'd12760: duty=167; 15'd12761: duty=173; 15'd12762: duty=174; 15'd12763: duty=170; 15'd12764: duty=170; 15'd12765: duty=163; 15'd12766: duty=159; 15'd12767: duty=156;
15'd12768: duty=156; 15'd12769: duty=159; 15'd12770: duty=151; 15'd12771: duty=152; 15'd12772: duty=156; 15'd12773: duty=151; 15'd12774: duty=140; 15'd12775: duty=137;
15'd12776: duty=137; 15'd12777: duty=142; 15'd12778: duty=139; 15'd12779: duty=136; 15'd12780: duty=133; 15'd12781: duty=124; 15'd12782: duty=126; 15'd12783: duty=119;
15'd12784: duty=110; 15'd12785: duty=119; 15'd12786: duty=115; 15'd12787: duty=109; 15'd12788: duty=112; 15'd12789: duty=107; 15'd12790: duty=101; 15'd12791: duty=93;
15'd12792: duty=90; 15'd12793: duty=91; 15'd12794: duty=86; 15'd12795: duty=88; 15'd12796: duty=90; 15'd12797: duty=90; 15'd12798: duty=87; 15'd12799: duty=91;
15'd12800: duty=90; 15'd12801: duty=85; 15'd12802: duty=96; 15'd12803: duty=101; 15'd12804: duty=110; 15'd12805: duty=110; 15'd12806: duty=99; 15'd12807: duty=98;
15'd12808: duty=98; 15'd12809: duty=107; 15'd12810: duty=115; 15'd12811: duty=114; 15'd12812: duty=115; 15'd12813: duty=116; 15'd12814: duty=112; 15'd12815: duty=114;
15'd12816: duty=118; 15'd12817: duty=117; 15'd12818: duty=119; 15'd12819: duty=116; 15'd12820: duty=116; 15'd12821: duty=121; 15'd12822: duty=119; 15'd12823: duty=121;
15'd12824: duty=136; 15'd12825: duty=139; 15'd12826: duty=147; 15'd12827: duty=143; 15'd12828: duty=147; 15'd12829: duty=149; 15'd12830: duty=142; 15'd12831: duty=153;
15'd12832: duty=142; 15'd12833: duty=145; 15'd12834: duty=148; 15'd12835: duty=149; 15'd12836: duty=151; 15'd12837: duty=153; 15'd12838: duty=148; 15'd12839: duty=156;
15'd12840: duty=161; 15'd12841: duty=157; 15'd12842: duty=162; 15'd12843: duty=162; 15'd12844: duty=165; 15'd12845: duty=153; 15'd12846: duty=156; 15'd12847: duty=167;
15'd12848: duty=165; 15'd12849: duty=168; 15'd12850: duty=173; 15'd12851: duty=163; 15'd12852: duty=161; 15'd12853: duty=165; 15'd12854: duty=163; 15'd12855: duty=159;
15'd12856: duty=162; 15'd12857: duty=161; 15'd12858: duty=156; 15'd12859: duty=151; 15'd12860: duty=149; 15'd12861: duty=150; 15'd12862: duty=151; 15'd12863: duty=156;
15'd12864: duty=153; 15'd12865: duty=147; 15'd12866: duty=148; 15'd12867: duty=141; 15'd12868: duty=131; 15'd12869: duty=127; 15'd12870: duty=120; 15'd12871: duty=121;
15'd12872: duty=122; 15'd12873: duty=121; 15'd12874: duty=121; 15'd12875: duty=113; 15'd12876: duty=113; 15'd12877: duty=110; 15'd12878: duty=104; 15'd12879: duty=98;
15'd12880: duty=94; 15'd12881: duty=95; 15'd12882: duty=96; 15'd12883: duty=96; 15'd12884: duty=91; 15'd12885: duty=95; 15'd12886: duty=95; 15'd12887: duty=101;
15'd12888: duty=102; 15'd12889: duty=93; 15'd12890: duty=101; 15'd12891: duty=104; 15'd12892: duty=104; 15'd12893: duty=104; 15'd12894: duty=99; 15'd12895: duty=98;
15'd12896: duty=96; 15'd12897: duty=102; 15'd12898: duty=110; 15'd12899: duty=114; 15'd12900: duty=115; 15'd12901: duty=104; 15'd12902: duty=105; 15'd12903: duty=102;
15'd12904: duty=99; 15'd12905: duty=107; 15'd12906: duty=109; 15'd12907: duty=113; 15'd12908: duty=118; 15'd12909: duty=122; 15'd12910: duty=124; 15'd12911: duty=128;
15'd12912: duty=128; 15'd12913: duty=133; 15'd12914: duty=126; 15'd12915: duty=129; 15'd12916: duty=134; 15'd12917: duty=127; 15'd12918: duty=134; 15'd12919: duty=132;
15'd12920: duty=139; 15'd12921: duty=146; 15'd12922: duty=142; 15'd12923: duty=146; 15'd12924: duty=154; 15'd12925: duty=165; 15'd12926: duty=171; 15'd12927: duty=163;
15'd12928: duty=164; 15'd12929: duty=171; 15'd12930: duty=161; 15'd12931: duty=168; 15'd12932: duty=168; 15'd12933: duty=157; 15'd12934: duty=159; 15'd12935: duty=157;
15'd12936: duty=171; 15'd12937: duty=171; 15'd12938: duty=164; 15'd12939: duty=164; 15'd12940: duty=163; 15'd12941: duty=163; 15'd12942: duty=166; 15'd12943: duty=162;
15'd12944: duty=159; 15'd12945: duty=154; 15'd12946: duty=154; 15'd12947: duty=159; 15'd12948: duty=160; 15'd12949: duty=163; 15'd12950: duty=165; 15'd12951: duty=166;
15'd12952: duty=159; 15'd12953: duty=159; 15'd12954: duty=153; 15'd12955: duty=142; 15'd12956: duty=137; 15'd12957: duty=134; 15'd12958: duty=131; 15'd12959: duty=127;
15'd12960: duty=119; 15'd12961: duty=114; 15'd12962: duty=104; 15'd12963: duty=102; 15'd12964: duty=106; 15'd12965: duty=102; 15'd12966: duty=102; 15'd12967: duty=104;
15'd12968: duty=104; 15'd12969: duty=99; 15'd12970: duty=98; 15'd12971: duty=96; 15'd12972: duty=90; 15'd12973: duty=93; 15'd12974: duty=90; 15'd12975: duty=95;
15'd12976: duty=90; 15'd12977: duty=90; 15'd12978: duty=92; 15'd12979: duty=90; 15'd12980: duty=95; 15'd12981: duty=94; 15'd12982: duty=98; 15'd12983: duty=100;
15'd12984: duty=104; 15'd12985: duty=104; 15'd12986: duty=110; 15'd12987: duty=104; 15'd12988: duty=103; 15'd12989: duty=107; 15'd12990: duty=106; 15'd12991: duty=110;
15'd12992: duty=115; 15'd12993: duty=118; 15'd12994: duty=118; 15'd12995: duty=115; 15'd12996: duty=118; 15'd12997: duty=119; 15'd12998: duty=125; 15'd12999: duty=135;
15'd13000: duty=134; 15'd13001: duty=128; 15'd13002: duty=127; 15'd13003: duty=129; 15'd13004: duty=124; 15'd13005: duty=136; 15'd13006: duty=139; 15'd13007: duty=144;
15'd13008: duty=153; 15'd13009: duty=143; 15'd13010: duty=151; 15'd13011: duty=153; 15'd13012: duty=151; 15'd13013: duty=157; 15'd13014: duty=157; 15'd13015: duty=165;
15'd13016: duty=170; 15'd13017: duty=157; 15'd13018: duty=151; 15'd13019: duty=157; 15'd13020: duty=157; 15'd13021: duty=168; 15'd13022: duty=168; 15'd13023: duty=168;
15'd13024: duty=173; 15'd13025: duty=179; 15'd13026: duty=174; 15'd13027: duty=169; 15'd13028: duty=160; 15'd13029: duty=157; 15'd13030: duty=162; 15'd13031: duty=157;
15'd13032: duty=159; 15'd13033: duty=153; 15'd13034: duty=148; 15'd13035: duty=149; 15'd13036: duty=153; 15'd13037: duty=148; 15'd13038: duty=153; 15'd13039: duty=154;
15'd13040: duty=148; 15'd13041: duty=148; 15'd13042: duty=139; 15'd13043: duty=128; 15'd13044: duty=127; 15'd13045: duty=119; 15'd13046: duty=113; 15'd13047: duty=116;
15'd13048: duty=110; 15'd13049: duty=113; 15'd13050: duty=113; 15'd13051: duty=107; 15'd13052: duty=109; 15'd13053: duty=102; 15'd13054: duty=101; 15'd13055: duty=105;
15'd13056: duty=105; 15'd13057: duty=111; 15'd13058: duty=104; 15'd13059: duty=102; 15'd13060: duty=104; 15'd13061: duty=110; 15'd13062: duty=104; 15'd13063: duty=101;
15'd13064: duty=109; 15'd13065: duty=108; 15'd13066: duty=113; 15'd13067: duty=109; 15'd13068: duty=104; 15'd13069: duty=106; 15'd13070: duty=103; 15'd13071: duty=105;
15'd13072: duty=107; 15'd13073: duty=115; 15'd13074: duty=112; 15'd13075: duty=104; 15'd13076: duty=99; 15'd13077: duty=93; 15'd13078: duty=98; 15'd13079: duty=105;
15'd13080: duty=113; 15'd13081: duty=116; 15'd13082: duty=110; 15'd13083: duty=112; 15'd13084: duty=116; 15'd13085: duty=113; 15'd13086: duty=118; 15'd13087: duty=126;
15'd13088: duty=134; 15'd13089: duty=128; 15'd13090: duty=134; 15'd13091: duty=150; 15'd13092: duty=145; 15'd13093: duty=139; 15'd13094: duty=145; 15'd13095: duty=147;
15'd13096: duty=145; 15'd13097: duty=133; 15'd13098: duty=142; 15'd13099: duty=155; 15'd13100: duty=148; 15'd13101: duty=155; 15'd13102: duty=152; 15'd13103: duty=144;
15'd13104: duty=154; 15'd13105: duty=158; 15'd13106: duty=154; 15'd13107: duty=156; 15'd13108: duty=159; 15'd13109: duty=168; 15'd13110: duty=163; 15'd13111: duty=166;
15'd13112: duty=177; 15'd13113: duty=170; 15'd13114: duty=171; 15'd13115: duty=168; 15'd13116: duty=163; 15'd13117: duty=167; 15'd13118: duty=168; 15'd13119: duty=161;
15'd13120: duty=158; 15'd13121: duty=156; 15'd13122: duty=148; 15'd13123: duty=144; 15'd13124: duty=145; 15'd13125: duty=151; 15'd13126: duty=144; 15'd13127: duty=148;
15'd13128: duty=149; 15'd13129: duty=144; 15'd13130: duty=146; 15'd13131: duty=136; 15'd13132: duty=134; 15'd13133: duty=130; 15'd13134: duty=125; 15'd13135: duty=115;
15'd13136: duty=116; 15'd13137: duty=118; 15'd13138: duty=111; 15'd13139: duty=103; 15'd13140: duty=102; 15'd13141: duty=107; 15'd13142: duty=102; 15'd13143: duty=98;
15'd13144: duty=100; 15'd13145: duty=107; 15'd13146: duty=101; 15'd13147: duty=106; 15'd13148: duty=104; 15'd13149: duty=90; 15'd13150: duty=90; 15'd13151: duty=92;
15'd13152: duty=96; 15'd13153: duty=98; 15'd13154: duty=101; 15'd13155: duty=107; 15'd13156: duty=105; 15'd13157: duty=106; 15'd13158: duty=111; 15'd13159: duty=106;
15'd13160: duty=105; 15'd13161: duty=107; 15'd13162: duty=108; 15'd13163: duty=112; 15'd13164: duty=117; 15'd13165: duty=112; 15'd13166: duty=122; 15'd13167: duty=126;
15'd13168: duty=116; 15'd13169: duty=121; 15'd13170: duty=125; 15'd13171: duty=118; 15'd13172: duty=116; 15'd13173: duty=118; 15'd13174: duty=116; 15'd13175: duty=126;
15'd13176: duty=127; 15'd13177: duty=131; 15'd13178: duty=133; 15'd13179: duty=133; 15'd13180: duty=145; 15'd13181: duty=139; 15'd13182: duty=131; 15'd13183: duty=134;
15'd13184: duty=145; 15'd13185: duty=139; 15'd13186: duty=145; 15'd13187: duty=160; 15'd13188: duty=153; 15'd13189: duty=145; 15'd13190: duty=143; 15'd13191: duty=154;
15'd13192: duty=160; 15'd13193: duty=156; 15'd13194: duty=151; 15'd13195: duty=159; 15'd13196: duty=159; 15'd13197: duty=153; 15'd13198: duty=153; 15'd13199: duty=150;
15'd13200: duty=153; 15'd13201: duty=157; 15'd13202: duty=157; 15'd13203: duty=167; 15'd13204: duty=165; 15'd13205: duty=160; 15'd13206: duty=163; 15'd13207: duty=162;
15'd13208: duty=159; 15'd13209: duty=163; 15'd13210: duty=165; 15'd13211: duty=157; 15'd13212: duty=160; 15'd13213: duty=160; 15'd13214: duty=156; 15'd13215: duty=146;
15'd13216: duty=139; 15'd13217: duty=133; 15'd13218: duty=131; 15'd13219: duty=127; 15'd13220: duty=124; 15'd13221: duty=116; 15'd13222: duty=116; 15'd13223: duty=122;
15'd13224: duty=116; 15'd13225: duty=115; 15'd13226: duty=118; 15'd13227: duty=111; 15'd13228: duty=117; 15'd13229: duty=118; 15'd13230: duty=115; 15'd13231: duty=114;
15'd13232: duty=103; 15'd13233: duty=110; 15'd13234: duty=104; 15'd13235: duty=97; 15'd13236: duty=106; 15'd13237: duty=107; 15'd13238: duty=102; 15'd13239: duty=115;
15'd13240: duty=107; 15'd13241: duty=96; 15'd13242: duty=101; 15'd13243: duty=101; 15'd13244: duty=113; 15'd13245: duty=110; 15'd13246: duty=99; 15'd13247: duty=108;
15'd13248: duty=112; 15'd13249: duty=105; 15'd13250: duty=119; 15'd13251: duty=124; 15'd13252: duty=107; 15'd13253: duty=111; 15'd13254: duty=124; 15'd13255: duty=114;
15'd13256: duty=111; 15'd13257: duty=121; 15'd13258: duty=119; 15'd13259: duty=122; 15'd13260: duty=118; 15'd13261: duty=116; 15'd13262: duty=110; 15'd13263: duty=107;
15'd13264: duty=121; 15'd13265: duty=136; 15'd13266: duty=140; 15'd13267: duty=142; 15'd13268: duty=137; 15'd13269: duty=139; 15'd13270: duty=157; 15'd13271: duty=147;
15'd13272: duty=143; 15'd13273: duty=150; 15'd13274: duty=145; 15'd13275: duty=142; 15'd13276: duty=140; 15'd13277: duty=142; 15'd13278: duty=142; 15'd13279: duty=144;
15'd13280: duty=155; 15'd13281: duty=153; 15'd13282: duty=155; 15'd13283: duty=161; 15'd13284: duty=160; 15'd13285: duty=170; 15'd13286: duty=174; 15'd13287: duty=170;
15'd13288: duty=159; 15'd13289: duty=152; 15'd13290: duty=165; 15'd13291: duty=172; 15'd13292: duty=163; 15'd13293: duty=156; 15'd13294: duty=157; 15'd13295: duty=150;
15'd13296: duty=152; 15'd13297: duty=158; 15'd13298: duty=154; 15'd13299: duty=152; 15'd13300: duty=158; 15'd13301: duty=156; 15'd13302: duty=151; 15'd13303: duty=147;
15'd13304: duty=139; 15'd13305: duty=131; 15'd13306: duty=128; 15'd13307: duty=127; 15'd13308: duty=125; 15'd13309: duty=124; 15'd13310: duty=121; 15'd13311: duty=118;
15'd13312: duty=116; 15'd13313: duty=118; 15'd13314: duty=111; 15'd13315: duty=107; 15'd13316: duty=104; 15'd13317: duty=98; 15'd13318: duty=99; 15'd13319: duty=96;
15'd13320: duty=98; 15'd13321: duty=104; 15'd13322: duty=90; 15'd13323: duty=87; 15'd13324: duty=89; 15'd13325: duty=93; 15'd13326: duty=105; 15'd13327: duty=99;
15'd13328: duty=101; 15'd13329: duty=104; 15'd13330: duty=106; 15'd13331: duty=107; 15'd13332: duty=109; 15'd13333: duty=108; 15'd13334: duty=109; 15'd13335: duty=118;
15'd13336: duty=121; 15'd13337: duty=121; 15'd13338: duty=128; 15'd13339: duty=119; 15'd13340: duty=110; 15'd13341: duty=125; 15'd13342: duty=124; 15'd13343: duty=130;
15'd13344: duty=124; 15'd13345: duty=112; 15'd13346: duty=118; 15'd13347: duty=119; 15'd13348: duty=127; 15'd13349: duty=130; 15'd13350: duty=122; 15'd13351: duty=121;
15'd13352: duty=134; 15'd13353: duty=137; 15'd13354: duty=133; 15'd13355: duty=136; 15'd13356: duty=137; 15'd13357: duty=141; 15'd13358: duty=142; 15'd13359: duty=151;
15'd13360: duty=154; 15'd13361: duty=142; 15'd13362: duty=142; 15'd13363: duty=144; 15'd13364: duty=152; 15'd13365: duty=157; 15'd13366: duty=163; 15'd13367: duty=168;
15'd13368: duty=166; 15'd13369: duty=161; 15'd13370: duty=162; 15'd13371: duty=162; 15'd13372: duty=166; 15'd13373: duty=170; 15'd13374: duty=163; 15'd13375: duty=165;
15'd13376: duty=169; 15'd13377: duty=173; 15'd13378: duty=166; 15'd13379: duty=158; 15'd13380: duty=149; 15'd13381: duty=153; 15'd13382: duty=165; 15'd13383: duty=167;
15'd13384: duty=160; 15'd13385: duty=155; 15'd13386: duty=151; 15'd13387: duty=148; 15'd13388: duty=139; 15'd13389: duty=138; 15'd13390: duty=139; 15'd13391: duty=133;
15'd13392: duty=131; 15'd13393: duty=134; 15'd13394: duty=127; 15'd13395: duty=115; 15'd13396: duty=116; 15'd13397: duty=115; 15'd13398: duty=111; 15'd13399: duty=106;
15'd13400: duty=108; 15'd13401: duty=101; 15'd13402: duty=98; 15'd13403: duty=101; 15'd13404: duty=100; 15'd13405: duty=90; 15'd13406: duty=96; 15'd13407: duty=103;
15'd13408: duty=103; 15'd13409: duty=106; 15'd13410: duty=110; 15'd13411: duty=121; 15'd13412: duty=110; 15'd13413: duty=103; 15'd13414: duty=104; 15'd13415: duty=98;
15'd13416: duty=105; 15'd13417: duty=108; 15'd13418: duty=100; 15'd13419: duty=94; 15'd13420: duty=102; 15'd13421: duty=110; 15'd13422: duty=97; 15'd13423: duty=86;
15'd13424: duty=87; 15'd13425: duty=98; 15'd13426: duty=113; 15'd13427: duty=126; 15'd13428: duty=122; 15'd13429: duty=116; 15'd13430: duty=119; 15'd13431: duty=110;
15'd13432: duty=104; 15'd13433: duty=124; 15'd13434: duty=128; 15'd13435: duty=115; 15'd13436: duty=116; 15'd13437: duty=125; 15'd13438: duty=136; 15'd13439: duty=128;
15'd13440: duty=133; 15'd13441: duty=137; 15'd13442: duty=136; 15'd13443: duty=143; 15'd13444: duty=147; 15'd13445: duty=148; 15'd13446: duty=140; 15'd13447: duty=148;
15'd13448: duty=153; 15'd13449: duty=162; 15'd13450: duty=156; 15'd13451: duty=163; 15'd13452: duty=182; 15'd13453: duty=170; 15'd13454: duty=161; 15'd13455: duty=164;
15'd13456: duty=161; 15'd13457: duty=165; 15'd13458: duty=165; 15'd13459: duty=168; 15'd13460: duty=170; 15'd13461: duty=162; 15'd13462: duty=173; 15'd13463: duty=173;
15'd13464: duty=159; 15'd13465: duty=162; 15'd13466: duty=166; 15'd13467: duty=168; 15'd13468: duty=171; 15'd13469: duty=167; 15'd13470: duty=163; 15'd13471: duty=156;
15'd13472: duty=154; 15'd13473: duty=153; 15'd13474: duty=148; 15'd13475: duty=134; 15'd13476: duty=129; 15'd13477: duty=130; 15'd13478: duty=129; 15'd13479: duty=120;
15'd13480: duty=125; 15'd13481: duty=127; 15'd13482: duty=124; 15'd13483: duty=126; 15'd13484: duty=114; 15'd13485: duty=112; 15'd13486: duty=114; 15'd13487: duty=107;
15'd13488: duty=111; 15'd13489: duty=121; 15'd13490: duty=107; 15'd13491: duty=103; 15'd13492: duty=111; 15'd13493: duty=101; 15'd13494: duty=93; 15'd13495: duty=93;
15'd13496: duty=93; 15'd13497: duty=104; 15'd13498: duty=99; 15'd13499: duty=95; 15'd13500: duty=93; 15'd13501: duty=95; 15'd13502: duty=87; 15'd13503: duty=98;
15'd13504: duty=105; 15'd13505: duty=99; 15'd13506: duty=107; 15'd13507: duty=107; 15'd13508: duty=118; 15'd13509: duty=121; 15'd13510: duty=113; 15'd13511: duty=102;
15'd13512: duty=111; 15'd13513: duty=119; 15'd13514: duty=133; 15'd13515: duty=139; 15'd13516: duty=127; 15'd13517: duty=124; 15'd13518: duty=118; 15'd13519: duty=99;
15'd13520: duty=100; 15'd13521: duty=105; 15'd13522: duty=106; 15'd13523: duty=120; 15'd13524: duty=121; 15'd13525: duty=116; 15'd13526: duty=123; 15'd13527: duty=132;
15'd13528: duty=130; 15'd13529: duty=131; 15'd13530: duty=142; 15'd13531: duty=157; 15'd13532: duty=167; 15'd13533: duty=160; 15'd13534: duty=157; 15'd13535: duty=150;
15'd13536: duty=143; 15'd13537: duty=153; 15'd13538: duty=154; 15'd13539: duty=151; 15'd13540: duty=156; 15'd13541: duty=158; 15'd13542: duty=154; 15'd13543: duty=161;
15'd13544: duty=166; 15'd13545: duty=170; 15'd13546: duty=161; 15'd13547: duty=165; 15'd13548: duty=179; 15'd13549: duty=173; 15'd13550: duty=172; 15'd13551: duty=174;
15'd13552: duty=163; 15'd13553: duty=164; 15'd13554: duty=168; 15'd13555: duty=164; 15'd13556: duty=168; 15'd13557: duty=161; 15'd13558: duty=157; 15'd13559: duty=161;
15'd13560: duty=155; 15'd13561: duty=146; 15'd13562: duty=137; 15'd13563: duty=127; 15'd13564: duty=127; 15'd13565: duty=124; 15'd13566: duty=119; 15'd13567: duty=118;
15'd13568: duty=119; 15'd13569: duty=109; 15'd13570: duty=111; 15'd13571: duty=122; 15'd13572: duty=113; 15'd13573: duty=115; 15'd13574: duty=114; 15'd13575: duty=108;
15'd13576: duty=113; 15'd13577: duty=110; 15'd13578: duty=101; 15'd13579: duty=96; 15'd13580: duty=101; 15'd13581: duty=95; 15'd13582: duty=100; 15'd13583: duty=102;
15'd13584: duty=93; 15'd13585: duty=102; 15'd13586: duty=98; 15'd13587: duty=101; 15'd13588: duty=115; 15'd13589: duty=96; 15'd13590: duty=98; 15'd13591: duty=102;
15'd13592: duty=87; 15'd13593: duty=96; 15'd13594: duty=112; 15'd13595: duty=96; 15'd13596: duty=97; 15'd13597: duty=104; 15'd13598: duty=107; 15'd13599: duty=116;
15'd13600: duty=110; 15'd13601: duty=127; 15'd13602: duty=119; 15'd13603: duty=118; 15'd13604: duty=123; 15'd13605: duty=131; 15'd13606: duty=120; 15'd13607: duty=117;
15'd13608: duty=136; 15'd13609: duty=133; 15'd13610: duty=134; 15'd13611: duty=136; 15'd13612: duty=136; 15'd13613: duty=126; 15'd13614: duty=139; 15'd13615: duty=148;
15'd13616: duty=139; 15'd13617: duty=142; 15'd13618: duty=156; 15'd13619: duty=151; 15'd13620: duty=157; 15'd13621: duty=163; 15'd13622: duty=162; 15'd13623: duty=163;
15'd13624: duty=160; 15'd13625: duty=164; 15'd13626: duty=165; 15'd13627: duty=156; 15'd13628: duty=160; 15'd13629: duty=168; 15'd13630: duty=170; 15'd13631: duty=176;
15'd13632: duty=183; 15'd13633: duty=176; 15'd13634: duty=172; 15'd13635: duty=165; 15'd13636: duty=159; 15'd13637: duty=160; 15'd13638: duty=163; 15'd13639: duty=167;
15'd13640: duty=163; 15'd13641: duty=161; 15'd13642: duty=166; 15'd13643: duty=167; 15'd13644: duty=156; 15'd13645: duty=151; 15'd13646: duty=145; 15'd13647: duty=142;
15'd13648: duty=137; 15'd13649: duty=143; 15'd13650: duty=133; 15'd13651: duty=126; 15'd13652: duty=119; 15'd13653: duty=112; 15'd13654: duty=116; 15'd13655: duty=102;
15'd13656: duty=104; 15'd13657: duty=101; 15'd13658: duty=95; 15'd13659: duty=98; 15'd13660: duty=98; 15'd13661: duty=104; 15'd13662: duty=106; 15'd13663: duty=96;
15'd13664: duty=92; 15'd13665: duty=88; 15'd13666: duty=92; 15'd13667: duty=89; 15'd13668: duty=84; 15'd13669: duty=90; 15'd13670: duty=95; 15'd13671: duty=97;
15'd13672: duty=86; 15'd13673: duty=86; 15'd13674: duty=103; 15'd13675: duty=102; 15'd13676: duty=106; 15'd13677: duty=99; 15'd13678: duty=100; 15'd13679: duty=105;
15'd13680: duty=109; 15'd13681: duty=116; 15'd13682: duty=111; 15'd13683: duty=122; 15'd13684: duty=126; 15'd13685: duty=119; 15'd13686: duty=127; 15'd13687: duty=132;
15'd13688: duty=123; 15'd13689: duty=122; 15'd13690: duty=117; 15'd13691: duty=119; 15'd13692: duty=127; 15'd13693: duty=125; 15'd13694: duty=123; 15'd13695: duty=134;
15'd13696: duty=137; 15'd13697: duty=145; 15'd13698: duty=136; 15'd13699: duty=137; 15'd13700: duty=144; 15'd13701: duty=141; 15'd13702: duty=149; 15'd13703: duty=155;
15'd13704: duty=159; 15'd13705: duty=150; 15'd13706: duty=153; 15'd13707: duty=156; 15'd13708: duty=164; 15'd13709: duty=167; 15'd13710: duty=159; 15'd13711: duty=163;
15'd13712: duty=168; 15'd13713: duty=168; 15'd13714: duty=167; 15'd13715: duty=156; 15'd13716: duty=169; 15'd13717: duty=171; 15'd13718: duty=171; 15'd13719: duty=179;
15'd13720: duty=176; 15'd13721: duty=176; 15'd13722: duty=165; 15'd13723: duty=167; 15'd13724: duty=168; 15'd13725: duty=163; 15'd13726: duty=167; 15'd13727: duty=163;
15'd13728: duty=159; 15'd13729: duty=159; 15'd13730: duty=144; 15'd13731: duty=128; 15'd13732: duty=126; 15'd13733: duty=129; 15'd13734: duty=124; 15'd13735: duty=125;
15'd13736: duty=126; 15'd13737: duty=122; 15'd13738: duty=118; 15'd13739: duty=119; 15'd13740: duty=109; 15'd13741: duty=110; 15'd13742: duty=114; 15'd13743: duty=111;
15'd13744: duty=114; 15'd13745: duty=108; 15'd13746: duty=104; 15'd13747: duty=103; 15'd13748: duty=95; 15'd13749: duty=87; 15'd13750: duty=90; 15'd13751: duty=92;
15'd13752: duty=89; 15'd13753: duty=108; 15'd13754: duty=107; 15'd13755: duty=94; 15'd13756: duty=95; 15'd13757: duty=86; 15'd13758: duty=83; 15'd13759: duty=84;
15'd13760: duty=100; 15'd13761: duty=108; 15'd13762: duty=113; 15'd13763: duty=114; 15'd13764: duty=107; 15'd13765: duty=100; 15'd13766: duty=101; 15'd13767: duty=105;
15'd13768: duty=111; 15'd13769: duty=114; 15'd13770: duty=114; 15'd13771: duty=128; 15'd13772: duty=126; 15'd13773: duty=116; 15'd13774: duty=104; 15'd13775: duty=100;
15'd13776: duty=114; 15'd13777: duty=130; 15'd13778: duty=131; 15'd13779: duty=138; 15'd13780: duty=133; 15'd13781: duty=137; 15'd13782: duty=148; 15'd13783: duty=151;
15'd13784: duty=152; 15'd13785: duty=146; 15'd13786: duty=139; 15'd13787: duty=142; 15'd13788: duty=161; 15'd13789: duty=166; 15'd13790: duty=153; 15'd13791: duty=141;
15'd13792: duty=143; 15'd13793: duty=156; 15'd13794: duty=167; 15'd13795: duty=166; 15'd13796: duty=159; 15'd13797: duty=154; 15'd13798: duty=156; 15'd13799: duty=151;
15'd13800: duty=166; 15'd13801: duty=174; 15'd13802: duty=174; 15'd13803: duty=172; 15'd13804: duty=153; 15'd13805: duty=168; 15'd13806: duty=174; 15'd13807: duty=171;
15'd13808: duty=171; 15'd13809: duty=167; 15'd13810: duty=167; 15'd13811: duty=173; 15'd13812: duty=185; 15'd13813: duty=170; 15'd13814: duty=159; 15'd13815: duty=148;
15'd13816: duty=142; 15'd13817: duty=142; 15'd13818: duty=135; 15'd13819: duty=128; 15'd13820: duty=134; 15'd13821: duty=136; 15'd13822: duty=125; 15'd13823: duty=128;
15'd13824: duty=125; 15'd13825: duty=113; 15'd13826: duty=107; 15'd13827: duty=104; 15'd13828: duty=111; 15'd13829: duty=111; 15'd13830: duty=107; 15'd13831: duty=110;
15'd13832: duty=97; 15'd13833: duty=99; 15'd13834: duty=91; 15'd13835: duty=88; 15'd13836: duty=94; 15'd13837: duty=96; 15'd13838: duty=89; 15'd13839: duty=85;
15'd13840: duty=84; 15'd13841: duty=79; 15'd13842: duty=87; 15'd13843: duty=90; 15'd13844: duty=83; 15'd13845: duty=88; 15'd13846: duty=101; 15'd13847: duty=110;
15'd13848: duty=116; 15'd13849: duty=104; 15'd13850: duty=97; 15'd13851: duty=105; 15'd13852: duty=121; 15'd13853: duty=136; 15'd13854: duty=125; 15'd13855: duty=118;
15'd13856: duty=128; 15'd13857: duty=128; 15'd13858: duty=131; 15'd13859: duty=126; 15'd13860: duty=124; 15'd13861: duty=117; 15'd13862: duty=128; 15'd13863: duty=133;
15'd13864: duty=141; 15'd13865: duty=142; 15'd13866: duty=132; 15'd13867: duty=124; 15'd13868: duty=113; 15'd13869: duty=130; 15'd13870: duty=137; 15'd13871: duty=127;
15'd13872: duty=128; 15'd13873: duty=139; 15'd13874: duty=142; 15'd13875: duty=147; 15'd13876: duty=136; 15'd13877: duty=142; 15'd13878: duty=145; 15'd13879: duty=142;
15'd13880: duty=152; 15'd13881: duty=163; 15'd13882: duty=153; 15'd13883: duty=140; 15'd13884: duty=147; 15'd13885: duty=151; 15'd13886: duty=159; 15'd13887: duty=157;
15'd13888: duty=156; 15'd13889: duty=166; 15'd13890: duty=162; 15'd13891: duty=176; 15'd13892: duty=182; 15'd13893: duty=184; 15'd13894: duty=182; 15'd13895: duty=175;
15'd13896: duty=182; 15'd13897: duty=171; 15'd13898: duty=170; 15'd13899: duty=168; 15'd13900: duty=163; 15'd13901: duty=160; 15'd13902: duty=158; 15'd13903: duty=160;
15'd13904: duty=141; 15'd13905: duty=140; 15'd13906: duty=148; 15'd13907: duty=142; 15'd13908: duty=135; 15'd13909: duty=124; 15'd13910: duty=118; 15'd13911: duty=120;
15'd13912: duty=120; 15'd13913: duty=110; 15'd13914: duty=115; 15'd13915: duty=116; 15'd13916: duty=110; 15'd13917: duty=107; 15'd13918: duty=115; 15'd13919: duty=101;
15'd13920: duty=96; 15'd13921: duty=97; 15'd13922: duty=93; 15'd13923: duty=98; 15'd13924: duty=97; 15'd13925: duty=93; 15'd13926: duty=88; 15'd13927: duty=78;
15'd13928: duty=71; 15'd13929: duty=87; 15'd13930: duty=91; 15'd13931: duty=89; 15'd13932: duty=90; 15'd13933: duty=96; 15'd13934: duty=100; 15'd13935: duty=99;
15'd13936: duty=95; 15'd13937: duty=104; 15'd13938: duty=99; 15'd13939: duty=98; 15'd13940: duty=118; 15'd13941: duty=120; 15'd13942: duty=116; 15'd13943: duty=112;
15'd13944: duty=99; 15'd13945: duty=102; 15'd13946: duty=123; 15'd13947: duty=130; 15'd13948: duty=133; 15'd13949: duty=125; 15'd13950: duty=126; 15'd13951: duty=147;
15'd13952: duty=145; 15'd13953: duty=130; 15'd13954: duty=136; 15'd13955: duty=142; 15'd13956: duty=139; 15'd13957: duty=143; 15'd13958: duty=150; 15'd13959: duty=154;
15'd13960: duty=140; 15'd13961: duty=135; 15'd13962: duty=151; 15'd13963: duty=162; 15'd13964: duty=171; 15'd13965: duty=168; 15'd13966: duty=162; 15'd13967: duty=163;
15'd13968: duty=173; 15'd13969: duty=172; 15'd13970: duty=167; 15'd13971: duty=165; 15'd13972: duty=170; 15'd13973: duty=174; 15'd13974: duty=177; 15'd13975: duty=173;
15'd13976: duty=172; 15'd13977: duty=172; 15'd13978: duty=164; 15'd13979: duty=168; 15'd13980: duty=171; 15'd13981: duty=172; 15'd13982: duty=174; 15'd13983: duty=177;
15'd13984: duty=173; 15'd13985: duty=163; 15'd13986: duty=148; 15'd13987: duty=145; 15'd13988: duty=141; 15'd13989: duty=140; 15'd13990: duty=132; 15'd13991: duty=142;
15'd13992: duty=135; 15'd13993: duty=120; 15'd13994: duty=115; 15'd13995: duty=111; 15'd13996: duty=115; 15'd13997: duty=115; 15'd13998: duty=106; 15'd13999: duty=99;
15'd14000: duty=107; 15'd14001: duty=105; 15'd14002: duty=112; 15'd14003: duty=92; 15'd14004: duty=75; 15'd14005: duty=80; 15'd14006: duty=94; 15'd14007: duty=91;
15'd14008: duty=92; 15'd14009: duty=88; 15'd14010: duty=78; 15'd14011: duty=82; 15'd14012: duty=83; 15'd14013: duty=86; 15'd14014: duty=95; 15'd14015: duty=91;
15'd14016: duty=95; 15'd14017: duty=99; 15'd14018: duty=100; 15'd14019: duty=111; 15'd14020: duty=107; 15'd14021: duty=108; 15'd14022: duty=106; 15'd14023: duty=114;
15'd14024: duty=112; 15'd14025: duty=114; 15'd14026: duty=107; 15'd14027: duty=109; 15'd14028: duty=112; 15'd14029: duty=105; 15'd14030: duty=124; 15'd14031: duty=125;
15'd14032: duty=124; 15'd14033: duty=127; 15'd14034: duty=124; 15'd14035: duty=123; 15'd14036: duty=125; 15'd14037: duty=134; 15'd14038: duty=139; 15'd14039: duty=146;
15'd14040: duty=161; 15'd14041: duty=155; 15'd14042: duty=158; 15'd14043: duty=162; 15'd14044: duty=156; 15'd14045: duty=168; 15'd14046: duty=147; 15'd14047: duty=150;
15'd14048: duty=159; 15'd14049: duty=153; 15'd14050: duty=163; 15'd14051: duty=165; 15'd14052: duty=175; 15'd14053: duty=170; 15'd14054: duty=172; 15'd14055: duty=170;
15'd14056: duty=173; 15'd14057: duty=163; 15'd14058: duty=153; 15'd14059: duty=167; 15'd14060: duty=174; 15'd14061: duty=167; 15'd14062: duty=181; 15'd14063: duty=181;
15'd14064: duty=169; 15'd14065: duty=166; 15'd14066: duty=177; 15'd14067: duty=182; 15'd14068: duty=169; 15'd14069: duty=170; 15'd14070: duty=150; 15'd14071: duty=138;
15'd14072: duty=137; 15'd14073: duty=126; 15'd14074: duty=121; 15'd14075: duty=117; 15'd14076: duty=117; 15'd14077: duty=116; 15'd14078: duty=119; 15'd14079: duty=125;
15'd14080: duty=131; 15'd14081: duty=124; 15'd14082: duty=114; 15'd14083: duty=123; 15'd14084: duty=120; 15'd14085: duty=112; 15'd14086: duty=105; 15'd14087: duty=103;
15'd14088: duty=103; 15'd14089: duty=95; 15'd14090: duty=96; 15'd14091: duty=106; 15'd14092: duty=93; 15'd14093: duty=97; 15'd14094: duty=93; 15'd14095: duty=81;
15'd14096: duty=91; 15'd14097: duty=106; 15'd14098: duty=102; 15'd14099: duty=92; 15'd14100: duty=90; 15'd14101: duty=98; 15'd14102: duty=102; 15'd14103: duty=92;
15'd14104: duty=107; 15'd14105: duty=102; 15'd14106: duty=92; 15'd14107: duty=86; 15'd14108: duty=99; 15'd14109: duty=97; 15'd14110: duty=93; 15'd14111: duty=93;
15'd14112: duty=92; 15'd14113: duty=99; 15'd14114: duty=109; 15'd14115: duty=109; 15'd14116: duty=115; 15'd14117: duty=124; 15'd14118: duty=127; 15'd14119: duty=131;
15'd14120: duty=142; 15'd14121: duty=134; 15'd14122: duty=129; 15'd14123: duty=136; 15'd14124: duty=139; 15'd14125: duty=140; 15'd14126: duty=138; 15'd14127: duty=158;
15'd14128: duty=160; 15'd14129: duty=165; 15'd14130: duty=159; 15'd14131: duty=167; 15'd14132: duty=172; 15'd14133: duty=165; 15'd14134: duty=166; 15'd14135: duty=157;
15'd14136: duty=161; 15'd14137: duty=165; 15'd14138: duty=152; 15'd14139: duty=147; 15'd14140: duty=160; 15'd14141: duty=169; 15'd14142: duty=166; 15'd14143: duty=176;
15'd14144: duty=183; 15'd14145: duty=176; 15'd14146: duty=174; 15'd14147: duty=182; 15'd14148: duty=184; 15'd14149: duty=178; 15'd14150: duty=177; 15'd14151: duty=172;
15'd14152: duty=173; 15'd14153: duty=176; 15'd14154: duty=169; 15'd14155: duty=164; 15'd14156: duty=158; 15'd14157: duty=144; 15'd14158: duty=144; 15'd14159: duty=140;
15'd14160: duty=140; 15'd14161: duty=133; 15'd14162: duty=126; 15'd14163: duty=117; 15'd14164: duty=108; 15'd14165: duty=114; 15'd14166: duty=107; 15'd14167: duty=105;
15'd14168: duty=105; 15'd14169: duty=93; 15'd14170: duty=103; 15'd14171: duty=108; 15'd14172: duty=116; 15'd14173: duty=110; 15'd14174: duty=99; 15'd14175: duty=104;
15'd14176: duty=104; 15'd14177: duty=98; 15'd14178: duty=86; 15'd14179: duty=80; 15'd14180: duty=78; 15'd14181: duty=94; 15'd14182: duty=93; 15'd14183: duty=98;
15'd14184: duty=92; 15'd14185: duty=96; 15'd14186: duty=110; 15'd14187: duty=105; 15'd14188: duty=91; 15'd14189: duty=93; 15'd14190: duty=95; 15'd14191: duty=95;
15'd14192: duty=106; 15'd14193: duty=116; 15'd14194: duty=112; 15'd14195: duty=100; 15'd14196: duty=106; 15'd14197: duty=118; 15'd14198: duty=119; 15'd14199: duty=107;
15'd14200: duty=119; 15'd14201: duty=124; 15'd14202: duty=126; 15'd14203: duty=122; 15'd14204: duty=113; 15'd14205: duty=110; 15'd14206: duty=125; 15'd14207: duty=127;
15'd14208: duty=133; 15'd14209: duty=136; 15'd14210: duty=139; 15'd14211: duty=145; 15'd14212: duty=137; 15'd14213: duty=137; 15'd14214: duty=146; 15'd14215: duty=154;
15'd14216: duty=146; 15'd14217: duty=158; 15'd14218: duty=163; 15'd14219: duty=162; 15'd14220: duty=174; 15'd14221: duty=173; 15'd14222: duty=168; 15'd14223: duty=165;
15'd14224: duty=156; 15'd14225: duty=168; 15'd14226: duty=168; 15'd14227: duty=161; 15'd14228: duty=166; 15'd14229: duty=164; 15'd14230: duty=166; 15'd14231: duty=165;
15'd14232: duty=173; 15'd14233: duty=182; 15'd14234: duty=178; 15'd14235: duty=177; 15'd14236: duty=187; 15'd14237: duty=182; 15'd14238: duty=158; 15'd14239: duty=150;
15'd14240: duty=155; 15'd14241: duty=155; 15'd14242: duty=151; 15'd14243: duty=145; 15'd14244: duty=145; 15'd14245: duty=138; 15'd14246: duty=136; 15'd14247: duty=130;
15'd14248: duty=127; 15'd14249: duty=121; 15'd14250: duty=120; 15'd14251: duty=121; 15'd14252: duty=119; 15'd14253: duty=117; 15'd14254: duty=118; 15'd14255: duty=120;
15'd14256: duty=107; 15'd14257: duty=116; 15'd14258: duty=121; 15'd14259: duty=116; 15'd14260: duty=98; 15'd14261: duty=101; 15'd14262: duty=108; 15'd14263: duty=90;
15'd14264: duty=98; 15'd14265: duty=90; 15'd14266: duty=79; 15'd14267: duty=93; 15'd14268: duty=102; 15'd14269: duty=90; 15'd14270: duty=86; 15'd14271: duty=98;
15'd14272: duty=96; 15'd14273: duty=95; 15'd14274: duty=98; 15'd14275: duty=108; 15'd14276: duty=106; 15'd14277: duty=88; 15'd14278: duty=98; 15'd14279: duty=111;
15'd14280: duty=107; 15'd14281: duty=98; 15'd14282: duty=103; 15'd14283: duty=92; 15'd14284: duty=93; 15'd14285: duty=119; 15'd14286: duty=128; 15'd14287: duty=129;
15'd14288: duty=124; 15'd14289: duty=120; 15'd14290: duty=128; 15'd14291: duty=138; 15'd14292: duty=124; 15'd14293: duty=131; 15'd14294: duty=133; 15'd14295: duty=136;
15'd14296: duty=126; 15'd14297: duty=131; 15'd14298: duty=148; 15'd14299: duty=149; 15'd14300: duty=142; 15'd14301: duty=146; 15'd14302: duty=171; 15'd14303: duty=167;
15'd14304: duty=168; 15'd14305: duty=156; 15'd14306: duty=159; 15'd14307: duty=171; 15'd14308: duty=181; 15'd14309: duty=180; 15'd14310: duty=170; 15'd14311: duty=174;
15'd14312: duty=170; 15'd14313: duty=173; 15'd14314: duty=171; 15'd14315: duty=170; 15'd14316: duty=173; 15'd14317: duty=165; 15'd14318: duty=179; 15'd14319: duty=168;
15'd14320: duty=162; 15'd14321: duty=165; 15'd14322: duty=167; 15'd14323: duty=161; 15'd14324: duty=157; 15'd14325: duty=154; 15'd14326: duty=149; 15'd14327: duty=159;
15'd14328: duty=155; 15'd14329: duty=150; 15'd14330: duty=138; 15'd14331: duty=124; 15'd14332: duty=128; 15'd14333: duty=133; 15'd14334: duty=125; 15'd14335: duty=129;
15'd14336: duty=122; 15'd14337: duty=118; 15'd14338: duty=112; 15'd14339: duty=120; 15'd14340: duty=107; 15'd14341: duty=96; 15'd14342: duty=98; 15'd14343: duty=104;
15'd14344: duty=98; 15'd14345: duty=88; 15'd14346: duty=89; 15'd14347: duty=88; 15'd14348: duty=81; 15'd14349: duty=81; 15'd14350: duty=93; 15'd14351: duty=87;
15'd14352: duty=90; 15'd14353: duty=89; 15'd14354: duty=92; 15'd14355: duty=96; 15'd14356: duty=95; 15'd14357: duty=84; 15'd14358: duty=99; 15'd14359: duty=111;
15'd14360: duty=110; 15'd14361: duty=102; 15'd14362: duty=100; 15'd14363: duty=114; 15'd14364: duty=122; 15'd14365: duty=114; 15'd14366: duty=113; 15'd14367: duty=107;
15'd14368: duty=93; 15'd14369: duty=104; 15'd14370: duty=109; 15'd14371: duty=112; 15'd14372: duty=107; 15'd14373: duty=110; 15'd14374: duty=128; 15'd14375: duty=124;
15'd14376: duty=128; 15'd14377: duty=136; 15'd14378: duty=150; 15'd14379: duty=153; 15'd14380: duty=148; 15'd14381: duty=161; 15'd14382: duty=159; 15'd14383: duty=153;
15'd14384: duty=159; 15'd14385: duty=154; 15'd14386: duty=153; 15'd14387: duty=163; 15'd14388: duty=171; 15'd14389: duty=166; 15'd14390: duty=156; 15'd14391: duty=156;
15'd14392: duty=154; 15'd14393: duty=156; 15'd14394: duty=158; 15'd14395: duty=166; 15'd14396: duty=171; 15'd14397: duty=169; 15'd14398: duty=175; 15'd14399: duty=177;
15'd14400: duty=169; 15'd14401: duty=177; 15'd14402: duty=181; 15'd14403: duty=184; 15'd14404: duty=173; 15'd14405: duty=163; 15'd14406: duty=176; 15'd14407: duty=167;
15'd14408: duty=155; 15'd14409: duty=149; 15'd14410: duty=144; 15'd14411: duty=140; 15'd14412: duty=130; 15'd14413: duty=127; 15'd14414: duty=120; 15'd14415: duty=116;
15'd14416: duty=126; 15'd14417: duty=123; 15'd14418: duty=121; 15'd14419: duty=125; 15'd14420: duty=115; 15'd14421: duty=115; 15'd14422: duty=121; 15'd14423: duty=116;
15'd14424: duty=106; 15'd14425: duty=101; 15'd14426: duty=107; 15'd14427: duty=105; 15'd14428: duty=101; 15'd14429: duty=86; 15'd14430: duty=91; 15'd14431: duty=101;
15'd14432: duty=102; 15'd14433: duty=112; 15'd14434: duty=99; 15'd14435: duty=93; 15'd14436: duty=93; 15'd14437: duty=95; 15'd14438: duty=105; 15'd14439: duty=107;
15'd14440: duty=111; 15'd14441: duty=120; 15'd14442: duty=117; 15'd14443: duty=109; 15'd14444: duty=108; 15'd14445: duty=106; 15'd14446: duty=100; 15'd14447: duty=98;
15'd14448: duty=110; 15'd14449: duty=113; 15'd14450: duty=122; 15'd14451: duty=117; 15'd14452: duty=111; 15'd14453: duty=118; 15'd14454: duty=125; 15'd14455: duty=124;
15'd14456: duty=124; 15'd14457: duty=136; 15'd14458: duty=116; 15'd14459: duty=113; 15'd14460: duty=125; 15'd14461: duty=126; 15'd14462: duty=132; 15'd14463: duty=133;
15'd14464: duty=121; 15'd14465: duty=136; 15'd14466: duty=141; 15'd14467: duty=139; 15'd14468: duty=154; 15'd14469: duty=168; 15'd14470: duty=167; 15'd14471: duty=162;
15'd14472: duty=159; 15'd14473: duty=156; 15'd14474: duty=164; 15'd14475: duty=157; 15'd14476: duty=147; 15'd14477: duty=154; 15'd14478: duty=153; 15'd14479: duty=157;
15'd14480: duty=170; 15'd14481: duty=166; 15'd14482: duty=170; 15'd14483: duty=165; 15'd14484: duty=173; 15'd14485: duty=171; 15'd14486: duty=164; 15'd14487: duty=171;
15'd14488: duty=167; 15'd14489: duty=169; 15'd14490: duty=173; 15'd14491: duty=172; 15'd14492: duty=170; 15'd14493: duty=155; 15'd14494: duty=150; 15'd14495: duty=149;
15'd14496: duty=147; 15'd14497: duty=141; 15'd14498: duty=130; 15'd14499: duty=128; 15'd14500: duty=127; 15'd14501: duty=125; 15'd14502: duty=120; 15'd14503: duty=116;
15'd14504: duty=98; 15'd14505: duty=114; 15'd14506: duty=118; 15'd14507: duty=112; 15'd14508: duty=107; 15'd14509: duty=112; 15'd14510: duty=112; 15'd14511: duty=117;
15'd14512: duty=120; 15'd14513: duty=105; 15'd14514: duty=101; 15'd14515: duty=99; 15'd14516: duty=107; 15'd14517: duty=104; 15'd14518: duty=100; 15'd14519: duty=101;
15'd14520: duty=95; 15'd14521: duty=87; 15'd14522: duty=76; 15'd14523: duty=88; 15'd14524: duty=103; 15'd14525: duty=98; 15'd14526: duty=106; 15'd14527: duty=96;
15'd14528: duty=89; 15'd14529: duty=98; 15'd14530: duty=112; 15'd14531: duty=124; 15'd14532: duty=113; 15'd14533: duty=102; 15'd14534: duty=116; 15'd14535: duty=125;
15'd14536: duty=127; 15'd14537: duty=112; 15'd14538: duty=113; 15'd14539: duty=124; 15'd14540: duty=125; 15'd14541: duty=118; 15'd14542: duty=113; 15'd14543: duty=123;
15'd14544: duty=128; 15'd14545: duty=119; 15'd14546: duty=128; 15'd14547: duty=134; 15'd14548: duty=132; 15'd14549: duty=139; 15'd14550: duty=134; 15'd14551: duty=147;
15'd14552: duty=145; 15'd14553: duty=139; 15'd14554: duty=143; 15'd14555: duty=148; 15'd14556: duty=148; 15'd14557: duty=155; 15'd14558: duty=159; 15'd14559: duty=155;
15'd14560: duty=162; 15'd14561: duty=161; 15'd14562: duty=162; 15'd14563: duty=168; 15'd14564: duty=165; 15'd14565: duty=185; 15'd14566: duty=179; 15'd14567: duty=175;
15'd14568: duty=172; 15'd14569: duty=176; 15'd14570: duty=180; 15'd14571: duty=164; 15'd14572: duty=180; 15'd14573: duty=169; 15'd14574: duty=166; 15'd14575: duty=172;
15'd14576: duty=165; 15'd14577: duty=159; 15'd14578: duty=152; 15'd14579: duty=141; 15'd14580: duty=155; 15'd14581: duty=157; 15'd14582: duty=149; 15'd14583: duty=140;
15'd14584: duty=129; 15'd14585: duty=133; 15'd14586: duty=122; 15'd14587: duty=118; 15'd14588: duty=118; 15'd14589: duty=124; 15'd14590: duty=116; 15'd14591: duty=114;
15'd14592: duty=119; 15'd14593: duty=118; 15'd14594: duty=112; 15'd14595: duty=113; 15'd14596: duty=106; 15'd14597: duty=98; 15'd14598: duty=100; 15'd14599: duty=93;
15'd14600: duty=104; 15'd14601: duty=102; 15'd14602: duty=87; 15'd14603: duty=81; 15'd14604: duty=92; 15'd14605: duty=87; 15'd14606: duty=89; 15'd14607: duty=91;
15'd14608: duty=94; 15'd14609: duty=108; 15'd14610: duty=107; 15'd14611: duty=105; 15'd14612: duty=107; 15'd14613: duty=103; 15'd14614: duty=94; 15'd14615: duty=96;
15'd14616: duty=106; 15'd14617: duty=98; 15'd14618: duty=101; 15'd14619: duty=110; 15'd14620: duty=97; 15'd14621: duty=102; 15'd14622: duty=104; 15'd14623: duty=114;
15'd14624: duty=121; 15'd14625: duty=126; 15'd14626: duty=126; 15'd14627: duty=125; 15'd14628: duty=133; 15'd14629: duty=129; 15'd14630: duty=127; 15'd14631: duty=127;
15'd14632: duty=120; 15'd14633: duty=138; 15'd14634: duty=141; 15'd14635: duty=138; 15'd14636: duty=155; 15'd14637: duty=140; 15'd14638: duty=135; 15'd14639: duty=154;
15'd14640: duty=153; 15'd14641: duty=148; 15'd14642: duty=148; 15'd14643: duty=158; 15'd14644: duty=171; 15'd14645: duty=162; 15'd14646: duty=161; 15'd14647: duty=165;
15'd14648: duty=173; 15'd14649: duty=177; 15'd14650: duty=187; 15'd14651: duty=177; 15'd14652: duty=167; 15'd14653: duty=171; 15'd14654: duty=174; 15'd14655: duty=169;
15'd14656: duty=161; 15'd14657: duty=157; 15'd14658: duty=164; 15'd14659: duty=165; 15'd14660: duty=159; 15'd14661: duty=163; 15'd14662: duty=168; 15'd14663: duty=168;
15'd14664: duty=162; 15'd14665: duty=160; 15'd14666: duty=150; 15'd14667: duty=149; 15'd14668: duty=147; 15'd14669: duty=145; 15'd14670: duty=133; 15'd14671: duty=128;
15'd14672: duty=124; 15'd14673: duty=124; 15'd14674: duty=130; 15'd14675: duty=130; 15'd14676: duty=121; 15'd14677: duty=127; 15'd14678: duty=115; 15'd14679: duty=107;
15'd14680: duty=108; 15'd14681: duty=99; 15'd14682: duty=91; 15'd14683: duty=95; 15'd14684: duty=94; 15'd14685: duty=93; 15'd14686: duty=97; 15'd14687: duty=92;
15'd14688: duty=96; 15'd14689: duty=96; 15'd14690: duty=102; 15'd14691: duty=84; 15'd14692: duty=96; 15'd14693: duty=77; 15'd14694: duty=85; 15'd14695: duty=92;
15'd14696: duty=77; 15'd14697: duty=84; 15'd14698: duty=83; 15'd14699: duty=95; 15'd14700: duty=100; 15'd14701: duty=117; 15'd14702: duty=124; 15'd14703: duty=123;
15'd14704: duty=119; 15'd14705: duty=123; 15'd14706: duty=125; 15'd14707: duty=124; 15'd14708: duty=119; 15'd14709: duty=110; 15'd14710: duty=113; 15'd14711: duty=103;
15'd14712: duty=114; 15'd14713: duty=127; 15'd14714: duty=134; 15'd14715: duty=135; 15'd14716: duty=128; 15'd14717: duty=132; 15'd14718: duty=146; 15'd14719: duty=150;
15'd14720: duty=148; 15'd14721: duty=151; 15'd14722: duty=142; 15'd14723: duty=150; 15'd14724: duty=148; 15'd14725: duty=156; 15'd14726: duty=145; 15'd14727: duty=159;
15'd14728: duty=154; 15'd14729: duty=154; 15'd14730: duty=171; 15'd14731: duty=171; 15'd14732: duty=179; 15'd14733: duty=170; 15'd14734: duty=168; 15'd14735: duty=163;
15'd14736: duty=153; 15'd14737: duty=165; 15'd14738: duty=163; 15'd14739: duty=149; 15'd14740: duty=161; 15'd14741: duty=166; 15'd14742: duty=178; 15'd14743: duty=186;
15'd14744: duty=178; 15'd14745: duty=174; 15'd14746: duty=174; 15'd14747: duty=174; 15'd14748: duty=173; 15'd14749: duty=163; 15'd14750: duty=161; 15'd14751: duty=144;
15'd14752: duty=139; 15'd14753: duty=141; 15'd14754: duty=131; 15'd14755: duty=122; 15'd14756: duty=116; 15'd14757: duty=111; 15'd14758: duty=121; 15'd14759: duty=116;
15'd14760: duty=109; 15'd14761: duty=97; 15'd14762: duty=97; 15'd14763: duty=97; 15'd14764: duty=97; 15'd14765: duty=111; 15'd14766: duty=104; 15'd14767: duty=110;
15'd14768: duty=117; 15'd14769: duty=108; 15'd14770: duty=106; 15'd14771: duty=97; 15'd14772: duty=86; 15'd14773: duty=91; 15'd14774: duty=95; 15'd14775: duty=94;
15'd14776: duty=90; 15'd14777: duty=91; 15'd14778: duty=81; 15'd14779: duty=101; 15'd14780: duty=106; 15'd14781: duty=94; 15'd14782: duty=97; 15'd14783: duty=111;
15'd14784: duty=117; 15'd14785: duty=110; 15'd14786: duty=97; 15'd14787: duty=105; 15'd14788: duty=109; 15'd14789: duty=111; 15'd14790: duty=115; 15'd14791: duty=122;
15'd14792: duty=130; 15'd14793: duty=129; 15'd14794: duty=120; 15'd14795: duty=118; 15'd14796: duty=118; 15'd14797: duty=114; 15'd14798: duty=127; 15'd14799: duty=113;
15'd14800: duty=124; 15'd14801: duty=128; 15'd14802: duty=129; 15'd14803: duty=155; 15'd14804: duty=154; 15'd14805: duty=146; 15'd14806: duty=145; 15'd14807: duty=143;
15'd14808: duty=156; 15'd14809: duty=150; 15'd14810: duty=158; 15'd14811: duty=172; 15'd14812: duty=162; 15'd14813: duty=166; 15'd14814: duty=171; 15'd14815: duty=168;
15'd14816: duty=162; 15'd14817: duty=154; 15'd14818: duty=153; 15'd14819: duty=163; 15'd14820: duty=165; 15'd14821: duty=166; 15'd14822: duty=164; 15'd14823: duty=158;
15'd14824: duty=173; 15'd14825: duty=177; 15'd14826: duty=162; 15'd14827: duty=162; 15'd14828: duty=179; 15'd14829: duty=180; 15'd14830: duty=172; 15'd14831: duty=172;
15'd14832: duty=159; 15'd14833: duty=160; 15'd14834: duty=171; 15'd14835: duty=169; 15'd14836: duty=158; 15'd14837: duty=157; 15'd14838: duty=148; 15'd14839: duty=132;
15'd14840: duty=124; 15'd14841: duty=114; 15'd14842: duty=109; 15'd14843: duty=105; 15'd14844: duty=100; 15'd14845: duty=103; 15'd14846: duty=102; 15'd14847: duty=102;
15'd14848: duty=97; 15'd14849: duty=95; 15'd14850: duty=89; 15'd14851: duty=97; 15'd14852: duty=100; 15'd14853: duty=88; 15'd14854: duty=97; 15'd14855: duty=100;
15'd14856: duty=95; 15'd14857: duty=91; 15'd14858: duty=91; 15'd14859: duty=86; 15'd14860: duty=91; 15'd14861: duty=83; 15'd14862: duty=92; 15'd14863: duty=103;
15'd14864: duty=108; 15'd14865: duty=109; 15'd14866: duty=123; 15'd14867: duty=112; 15'd14868: duty=83; 15'd14869: duty=91; 15'd14870: duty=94; 15'd14871: duty=92;
15'd14872: duty=109; 15'd14873: duty=117; 15'd14874: duty=115; 15'd14875: duty=125; 15'd14876: duty=125; 15'd14877: duty=123; 15'd14878: duty=125; 15'd14879: duty=135;
15'd14880: duty=132; 15'd14881: duty=129; 15'd14882: duty=130; 15'd14883: duty=141; 15'd14884: duty=136; 15'd14885: duty=139; 15'd14886: duty=143; 15'd14887: duty=137;
15'd14888: duty=130; 15'd14889: duty=126; 15'd14890: duty=128; 15'd14891: duty=129; 15'd14892: duty=135; 15'd14893: duty=146; 15'd14894: duty=147; 15'd14895: duty=142;
15'd14896: duty=138; 15'd14897: duty=147; 15'd14898: duty=150; 15'd14899: duty=151; 15'd14900: duty=158; 15'd14901: duty=169; 15'd14902: duty=172; 15'd14903: duty=168;
15'd14904: duty=173; 15'd14905: duty=162; 15'd14906: duty=169; 15'd14907: duty=165; 15'd14908: duty=169; 15'd14909: duty=160; 15'd14910: duty=164; 15'd14911: duty=174;
15'd14912: duty=167; 15'd14913: duty=171; 15'd14914: duty=168; 15'd14915: duty=163; 15'd14916: duty=163; 15'd14917: duty=163; 15'd14918: duty=170; 15'd14919: duty=168;
15'd14920: duty=150; 15'd14921: duty=155; 15'd14922: duty=156; 15'd14923: duty=144; 15'd14924: duty=144; 15'd14925: duty=132; 15'd14926: duty=132; 15'd14927: duty=134;
15'd14928: duty=118; 15'd14929: duty=120; 15'd14930: duty=121; 15'd14931: duty=124; 15'd14932: duty=111; 15'd14933: duty=111; 15'd14934: duty=109; 15'd14935: duty=99;
15'd14936: duty=109; 15'd14937: duty=99; 15'd14938: duty=100; 15'd14939: duty=90; 15'd14940: duty=76; 15'd14941: duty=87; 15'd14942: duty=89; 15'd14943: duty=91;
15'd14944: duty=84; 15'd14945: duty=87; 15'd14946: duty=87; 15'd14947: duty=88; 15'd14948: duty=98; 15'd14949: duty=97; 15'd14950: duty=98; 15'd14951: duty=108;
15'd14952: duty=104; 15'd14953: duty=99; 15'd14954: duty=101; 15'd14955: duty=102; 15'd14956: duty=110; 15'd14957: duty=105; 15'd14958: duty=100; 15'd14959: duty=102;
15'd14960: duty=109; 15'd14961: duty=114; 15'd14962: duty=107; 15'd14963: duty=116; 15'd14964: duty=131; 15'd14965: duty=127; 15'd14966: duty=126; 15'd14967: duty=127;
15'd14968: duty=116; 15'd14969: duty=119; 15'd14970: duty=130; 15'd14971: duty=139; 15'd14972: duty=142; 15'd14973: duty=137; 15'd14974: duty=142; 15'd14975: duty=151;
15'd14976: duty=145; 15'd14977: duty=151; 15'd14978: duty=163; 15'd14979: duty=150; 15'd14980: duty=146; 15'd14981: duty=143; 15'd14982: duty=147; 15'd14983: duty=154;
15'd14984: duty=140; 15'd14985: duty=149; 15'd14986: duty=162; 15'd14987: duty=163; 15'd14988: duty=174; 15'd14989: duty=166; 15'd14990: duty=171; 15'd14991: duty=169;
15'd14992: duty=165; 15'd14993: duty=184; 15'd14994: duty=177; 15'd14995: duty=176; 15'd14996: duty=177; 15'd14997: duty=169; 15'd14998: duty=179; 15'd14999: duty=172;
15'd15000: duty=161; 15'd15001: duty=160; 15'd15002: duty=165; 15'd15003: duty=168; 15'd15004: duty=170; 15'd15005: duty=168; 15'd15006: duty=153; 15'd15007: duty=157;
15'd15008: duty=165; 15'd15009: duty=162; 15'd15010: duty=145; 15'd15011: duty=139; 15'd15012: duty=126; 15'd15013: duty=128; 15'd15014: duty=136; 15'd15015: duty=116;
15'd15016: duty=115; 15'd15017: duty=111; 15'd15018: duty=113; 15'd15019: duty=110; 15'd15020: duty=107; 15'd15021: duty=108; 15'd15022: duty=100; 15'd15023: duty=95;
15'd15024: duty=86; 15'd15025: duty=87; 15'd15026: duty=87; 15'd15027: duty=82; 15'd15028: duty=81; 15'd15029: duty=85; 15'd15030: duty=76; 15'd15031: duty=79;
15'd15032: duty=75; 15'd15033: duty=82; 15'd15034: duty=90; 15'd15035: duty=85; 15'd15036: duty=99; 15'd15037: duty=105; 15'd15038: duty=98; 15'd15039: duty=101;
15'd15040: duty=104; 15'd15041: duty=96; 15'd15042: duty=104; 15'd15043: duty=105; 15'd15044: duty=116; 15'd15045: duty=107; 15'd15046: duty=116; 15'd15047: duty=127;
15'd15048: duty=116; 15'd15049: duty=112; 15'd15050: duty=113; 15'd15051: duty=121; 15'd15052: duty=125; 15'd15053: duty=123; 15'd15054: duty=124; 15'd15055: duty=123;
15'd15056: duty=124; 15'd15057: duty=139; 15'd15058: duty=124; 15'd15059: duty=126; 15'd15060: duty=134; 15'd15061: duty=133; 15'd15062: duty=138; 15'd15063: duty=142;
15'd15064: duty=145; 15'd15065: duty=136; 15'd15066: duty=138; 15'd15067: duty=155; 15'd15068: duty=168; 15'd15069: duty=166; 15'd15070: duty=157; 15'd15071: duty=172;
15'd15072: duty=165; 15'd15073: duty=159; 15'd15074: duty=174; 15'd15075: duty=170; 15'd15076: duty=168; 15'd15077: duty=169; 15'd15078: duty=168; 15'd15079: duty=167;
15'd15080: duty=165; 15'd15081: duty=170; 15'd15082: duty=175; 15'd15083: duty=167; 15'd15084: duty=172; 15'd15085: duty=177; 15'd15086: duty=178; 15'd15087: duty=176;
15'd15088: duty=182; 15'd15089: duty=190; 15'd15090: duty=183; 15'd15091: duty=176; 15'd15092: duty=176; 15'd15093: duty=164; 15'd15094: duty=151; 15'd15095: duty=154;
15'd15096: duty=143; 15'd15097: duty=137; 15'd15098: duty=125; 15'd15099: duty=113; 15'd15100: duty=124; 15'd15101: duty=129; 15'd15102: duty=112; 15'd15103: duty=112;
15'd15104: duty=114; 15'd15105: duty=113; 15'd15106: duty=112; 15'd15107: duty=107; 15'd15108: duty=110; 15'd15109: duty=96; 15'd15110: duty=98; 15'd15111: duty=99;
15'd15112: duty=90; 15'd15113: duty=98; 15'd15114: duty=87; 15'd15115: duty=84; 15'd15116: duty=98; 15'd15117: duty=82; 15'd15118: duty=85; 15'd15119: duty=91;
15'd15120: duty=104; 15'd15121: duty=102; 15'd15122: duty=84; 15'd15123: duty=100; 15'd15124: duty=98; 15'd15125: duty=90; 15'd15126: duty=84; 15'd15127: duty=78;
15'd15128: duty=85; 15'd15129: duty=98; 15'd15130: duty=105; 15'd15131: duty=113; 15'd15132: duty=104; 15'd15133: duty=98; 15'd15134: duty=107; 15'd15135: duty=106;
15'd15136: duty=110; 15'd15137: duty=115; 15'd15138: duty=123; 15'd15139: duty=121; 15'd15140: duty=116; 15'd15141: duty=123; 15'd15142: duty=128; 15'd15143: duty=126;
15'd15144: duty=128; 15'd15145: duty=138; 15'd15146: duty=137; 15'd15147: duty=138; 15'd15148: duty=141; 15'd15149: duty=142; 15'd15150: duty=146; 15'd15151: duty=148;
15'd15152: duty=149; 15'd15153: duty=146; 15'd15154: duty=160; 15'd15155: duty=162; 15'd15156: duty=158; 15'd15157: duty=161; 15'd15158: duty=163; 15'd15159: duty=169;
15'd15160: duty=169; 15'd15161: duty=169; 15'd15162: duty=160; 15'd15163: duty=169; 15'd15164: duty=177; 15'd15165: duty=167; 15'd15166: duty=173; 15'd15167: duty=176;
15'd15168: duty=171; 15'd15169: duty=162; 15'd15170: duty=174; 15'd15171: duty=179; 15'd15172: duty=174; 15'd15173: duty=173; 15'd15174: duty=165; 15'd15175: duty=173;
15'd15176: duty=176; 15'd15177: duty=169; 15'd15178: duty=165; 15'd15179: duty=157; 15'd15180: duty=148; 15'd15181: duty=148; 15'd15182: duty=143; 15'd15183: duty=134;
15'd15184: duty=134; 15'd15185: duty=128; 15'd15186: duty=119; 15'd15187: duty=121; 15'd15188: duty=122; 15'd15189: duty=124; 15'd15190: duty=116; 15'd15191: duty=113;
15'd15192: duty=118; 15'd15193: duty=118; 15'd15194: duty=110; 15'd15195: duty=100; 15'd15196: duty=102; 15'd15197: duty=98; 15'd15198: duty=94; 15'd15199: duty=95;
15'd15200: duty=93; 15'd15201: duty=84; 15'd15202: duty=85; 15'd15203: duty=74; 15'd15204: duty=83; 15'd15205: duty=84; 15'd15206: duty=83; 15'd15207: duty=100;
15'd15208: duty=92; 15'd15209: duty=106; 15'd15210: duty=98; 15'd15211: duty=89; 15'd15212: duty=92; 15'd15213: duty=89; 15'd15214: duty=95; 15'd15215: duty=105;
15'd15216: duty=106; 15'd15217: duty=100; 15'd15218: duty=99; 15'd15219: duty=111; 15'd15220: duty=119; 15'd15221: duty=124; 15'd15222: duty=120; 15'd15223: duty=117;
15'd15224: duty=120; 15'd15225: duty=118; 15'd15226: duty=128; 15'd15227: duty=135; 15'd15228: duty=137; 15'd15229: duty=126; 15'd15230: duty=142; 15'd15231: duty=142;
15'd15232: duty=136; 15'd15233: duty=133; 15'd15234: duty=130; 15'd15235: duty=140; 15'd15236: duty=144; 15'd15237: duty=143; 15'd15238: duty=147; 15'd15239: duty=148;
15'd15240: duty=136; 15'd15241: duty=143; 15'd15242: duty=153; 15'd15243: duty=151; 15'd15244: duty=158; 15'd15245: duty=154; 15'd15246: duty=157; 15'd15247: duty=177;
15'd15248: duty=187; 15'd15249: duty=186; 15'd15250: duty=168; 15'd15251: duty=161; 15'd15252: duty=173; 15'd15253: duty=179; 15'd15254: duty=181; 15'd15255: duty=179;
15'd15256: duty=178; 15'd15257: duty=175; 15'd15258: duty=168; 15'd15259: duty=173; 15'd15260: duty=164; 15'd15261: duty=157; 15'd15262: duty=156; 15'd15263: duty=151;
15'd15264: duty=145; 15'd15265: duty=156; 15'd15266: duty=154; 15'd15267: duty=143; 15'd15268: duty=142; 15'd15269: duty=133; 15'd15270: duty=133; 15'd15271: duty=131;
15'd15272: duty=130; 15'd15273: duty=133; 15'd15274: duty=132; 15'd15275: duty=123; 15'd15276: duty=124; 15'd15277: duty=117; 15'd15278: duty=108; 15'd15279: duty=107;
15'd15280: duty=108; 15'd15281: duty=92; 15'd15282: duty=98; 15'd15283: duty=98; 15'd15284: duty=93; 15'd15285: duty=106; 15'd15286: duty=86; 15'd15287: duty=86;
15'd15288: duty=96; 15'd15289: duty=112; 15'd15290: duty=114; 15'd15291: duty=101; 15'd15292: duty=94; 15'd15293: duty=95; 15'd15294: duty=85; 15'd15295: duty=81;
15'd15296: duty=81; 15'd15297: duty=83; 15'd15298: duty=88; 15'd15299: duty=89; 15'd15300: duty=95; 15'd15301: duty=111; 15'd15302: duty=119; 15'd15303: duty=110;
15'd15304: duty=114; 15'd15305: duty=112; 15'd15306: duty=112; 15'd15307: duty=115; 15'd15308: duty=118; 15'd15309: duty=114; 15'd15310: duty=119; 15'd15311: duty=112;
15'd15312: duty=110; 15'd15313: duty=110; 15'd15314: duty=118; 15'd15315: duty=124; 15'd15316: duty=139; 15'd15317: duty=150; 15'd15318: duty=138; 15'd15319: duty=133;
15'd15320: duty=136; 15'd15321: duty=144; 15'd15322: duty=142; 15'd15323: duty=151; 15'd15324: duty=154; 15'd15325: duty=164; 15'd15326: duty=165; 15'd15327: duty=157;
15'd15328: duty=157; 15'd15329: duty=164; 15'd15330: duty=154; 15'd15331: duty=162; 15'd15332: duty=171; 15'd15333: duty=173; 15'd15334: duty=173; 15'd15335: duty=167;
15'd15336: duty=167; 15'd15337: duty=161; 15'd15338: duty=160; 15'd15339: duty=167; 15'd15340: duty=175; 15'd15341: duty=175; 15'd15342: duty=174; 15'd15343: duty=168;
15'd15344: duty=169; 15'd15345: duty=165; 15'd15346: duty=175; 15'd15347: duty=178; 15'd15348: duty=173; 15'd15349: duty=166; 15'd15350: duty=163; 15'd15351: duty=159;
15'd15352: duty=152; 15'd15353: duty=142; 15'd15354: duty=142; 15'd15355: duty=136; 15'd15356: duty=127; 15'd15357: duty=127; 15'd15358: duty=124; 15'd15359: duty=127;
15'd15360: duty=121; 15'd15361: duty=115; 15'd15362: duty=108; 15'd15363: duty=101; 15'd15364: duty=104; 15'd15365: duty=102; 15'd15366: duty=93; 15'd15367: duty=108;
15'd15368: duty=105; 15'd15369: duty=81; 15'd15370: duty=90; 15'd15371: duty=99; 15'd15372: duty=95; 15'd15373: duty=93; 15'd15374: duty=87; 15'd15375: duty=91;
15'd15376: duty=90; 15'd15377: duty=96; 15'd15378: duty=81; 15'd15379: duty=63; 15'd15380: duty=81; 15'd15381: duty=90; 15'd15382: duty=101; 15'd15383: duty=113;
15'd15384: duty=102; 15'd15385: duty=109; 15'd15386: duty=121; 15'd15387: duty=114; 15'd15388: duty=117; 15'd15389: duty=119; 15'd15390: duty=111; 15'd15391: duty=113;
15'd15392: duty=129; 15'd15393: duty=111; 15'd15394: duty=103; 15'd15395: duty=114; 15'd15396: duty=112; 15'd15397: duty=112; 15'd15398: duty=119; 15'd15399: duty=126;
15'd15400: duty=126; 15'd15401: duty=132; 15'd15402: duty=138; 15'd15403: duty=142; 15'd15404: duty=154; 15'd15405: duty=142; 15'd15406: duty=146; 15'd15407: duty=147;
15'd15408: duty=143; 15'd15409: duty=159; 15'd15410: duty=160; 15'd15411: duty=160; 15'd15412: duty=157; 15'd15413: duty=163; 15'd15414: duty=175; 15'd15415: duty=172;
15'd15416: duty=170; 15'd15417: duty=164; 15'd15418: duty=162; 15'd15419: duty=172; 15'd15420: duty=167; 15'd15421: duty=169; 15'd15422: duty=165; 15'd15423: duty=162;
15'd15424: duty=169; 15'd15425: duty=169; 15'd15426: duty=178; 15'd15427: duty=188; 15'd15428: duty=176; 15'd15429: duty=174; 15'd15430: duty=174; 15'd15431: duty=168;
15'd15432: duty=170; 15'd15433: duty=164; 15'd15434: duty=150; 15'd15435: duty=136; 15'd15436: duty=128; 15'd15437: duty=122; 15'd15438: duty=131; 15'd15439: duty=122;
15'd15440: duty=116; 15'd15441: duty=126; 15'd15442: duty=129; 15'd15443: duty=123; 15'd15444: duty=116; 15'd15445: duty=119; 15'd15446: duty=119; 15'd15447: duty=107;
15'd15448: duty=111; 15'd15449: duty=116; 15'd15450: duty=123; 15'd15451: duty=110; 15'd15452: duty=96; 15'd15453: duty=93; 15'd15454: duty=91; 15'd15455: duty=101;
15'd15456: duty=95; 15'd15457: duty=84; 15'd15458: duty=103; 15'd15459: duty=105; 15'd15460: duty=102; 15'd15461: duty=101; 15'd15462: duty=92; 15'd15463: duty=98;
15'd15464: duty=96; 15'd15465: duty=107; 15'd15466: duty=100; 15'd15467: duty=93; 15'd15468: duty=86; 15'd15469: duty=88; 15'd15470: duty=103; 15'd15471: duty=104;
15'd15472: duty=109; 15'd15473: duty=107; 15'd15474: duty=103; 15'd15475: duty=114; 15'd15476: duty=112; 15'd15477: duty=105; 15'd15478: duty=103; 15'd15479: duty=105;
15'd15480: duty=115; 15'd15481: duty=108; 15'd15482: duty=109; 15'd15483: duty=127; 15'd15484: duty=133; 15'd15485: duty=129; 15'd15486: duty=121; 15'd15487: duty=132;
15'd15488: duty=137; 15'd15489: duty=141; 15'd15490: duty=158; 15'd15491: duty=152; 15'd15492: duty=147; 15'd15493: duty=146; 15'd15494: duty=154; 15'd15495: duty=151;
15'd15496: duty=157; 15'd15497: duty=169; 15'd15498: duty=165; 15'd15499: duty=168; 15'd15500: duty=162; 15'd15501: duty=174; 15'd15502: duty=178; 15'd15503: duty=175;
15'd15504: duty=175; 15'd15505: duty=176; 15'd15506: duty=180; 15'd15507: duty=182; 15'd15508: duty=180; 15'd15509: duty=168; 15'd15510: duty=166; 15'd15511: duty=170;
15'd15512: duty=171; 15'd15513: duty=174; 15'd15514: duty=177; 15'd15515: duty=176; 15'd15516: duty=176; 15'd15517: duty=170; 15'd15518: duty=165; 15'd15519: duty=158;
15'd15520: duty=154; 15'd15521: duty=153; 15'd15522: duty=148; 15'd15523: duty=139; 15'd15524: duty=135; 15'd15525: duty=137; 15'd15526: duty=132; 15'd15527: duty=123;
15'd15528: duty=126; 15'd15529: duty=125; 15'd15530: duty=114; 15'd15531: duty=111; 15'd15532: duty=108; 15'd15533: duty=113; 15'd15534: duty=105; 15'd15535: duty=98;
15'd15536: duty=95; 15'd15537: duty=90; 15'd15538: duty=87; 15'd15539: duty=93; 15'd15540: duty=88; 15'd15541: duty=94; 15'd15542: duty=87; 15'd15543: duty=89;
15'd15544: duty=99; 15'd15545: duty=97; 15'd15546: duty=102; 15'd15547: duty=93; 15'd15548: duty=86; 15'd15549: duty=87; 15'd15550: duty=89; 15'd15551: duty=82;
15'd15552: duty=89; 15'd15553: duty=90; 15'd15554: duty=95; 15'd15555: duty=104; 15'd15556: duty=114; 15'd15557: duty=103; 15'd15558: duty=109; 15'd15559: duty=113;
15'd15560: duty=111; 15'd15561: duty=99; 15'd15562: duty=97; 15'd15563: duty=110; 15'd15564: duty=111; 15'd15565: duty=117; 15'd15566: duty=124; 15'd15567: duty=135;
15'd15568: duty=137; 15'd15569: duty=132; 15'd15570: duty=134; 15'd15571: duty=135; 15'd15572: duty=121; 15'd15573: duty=122; 15'd15574: duty=128; 15'd15575: duty=129;
15'd15576: duty=120; 15'd15577: duty=138; 15'd15578: duty=151; 15'd15579: duty=137; 15'd15580: duty=142; 15'd15581: duty=144; 15'd15582: duty=150; 15'd15583: duty=160;
15'd15584: duty=155; 15'd15585: duty=166; 15'd15586: duty=173; 15'd15587: duty=175; 15'd15588: duty=182; 15'd15589: duty=172; 15'd15590: duty=161; 15'd15591: duty=171;
15'd15592: duty=176; 15'd15593: duty=179; 15'd15594: duty=191; 15'd15595: duty=182; 15'd15596: duty=187; 15'd15597: duty=191; 15'd15598: duty=174; 15'd15599: duty=171;
15'd15600: duty=174; 15'd15601: duty=177; 15'd15602: duty=165; 15'd15603: duty=160; 15'd15604: duty=159; 15'd15605: duty=153; 15'd15606: duty=142; 15'd15607: duty=133;
15'd15608: duty=137; 15'd15609: duty=133; 15'd15610: duty=133; 15'd15611: duty=135; 15'd15612: duty=139; 15'd15613: duty=124; 15'd15614: duty=128; 15'd15615: duty=130;
15'd15616: duty=127; 15'd15617: duty=123; 15'd15618: duty=114; 15'd15619: duty=117; 15'd15620: duty=110; 15'd15621: duty=105; 15'd15622: duty=114; 15'd15623: duty=107;
15'd15624: duty=93; 15'd15625: duty=90; 15'd15626: duty=91; 15'd15627: duty=101; 15'd15628: duty=110; 15'd15629: duty=98; 15'd15630: duty=84; 15'd15631: duty=88;
15'd15632: duty=79; 15'd15633: duty=73; 15'd15634: duty=77; 15'd15635: duty=81; 15'd15636: duty=99; 15'd15637: duty=118; 15'd15638: duty=104; 15'd15639: duty=106;
15'd15640: duty=111; 15'd15641: duty=107; 15'd15642: duty=113; 15'd15643: duty=116; 15'd15644: duty=126; 15'd15645: duty=106; 15'd15646: duty=90; 15'd15647: duty=79;
15'd15648: duty=81; 15'd15649: duty=107; 15'd15650: duty=107; 15'd15651: duty=113; 15'd15652: duty=119; 15'd15653: duty=128; 15'd15654: duty=131; 15'd15655: duty=144;
15'd15656: duty=142; 15'd15657: duty=127; 15'd15658: duty=143; 15'd15659: duty=147; 15'd15660: duty=150; 15'd15661: duty=157; 15'd15662: duty=150; 15'd15663: duty=141;
15'd15664: duty=136; 15'd15665: duty=145; 15'd15666: duty=159; 15'd15667: duty=162; 15'd15668: duty=157; 15'd15669: duty=148; 15'd15670: duty=150; 15'd15671: duty=158;
15'd15672: duty=161; 15'd15673: duty=154; 15'd15674: duty=159; 15'd15675: duty=174; 15'd15676: duty=165; 15'd15677: duty=165; 15'd15678: duty=182; 15'd15679: duty=181;
15'd15680: duty=176; 15'd15681: duty=172; 15'd15682: duty=181; 15'd15683: duty=186; 15'd15684: duty=184; 15'd15685: duty=189; 15'd15686: duty=181; 15'd15687: duty=175;
15'd15688: duty=168; 15'd15689: duty=158; 15'd15690: duty=151; 15'd15691: duty=143; 15'd15692: duty=140; 15'd15693: duty=140; 15'd15694: duty=145; 15'd15695: duty=137;
15'd15696: duty=138; 15'd15697: duty=129; 15'd15698: duty=116; 15'd15699: duty=119; 15'd15700: duty=124; 15'd15701: duty=124; 15'd15702: duty=123; 15'd15703: duty=121;
15'd15704: duty=114; 15'd15705: duty=117; 15'd15706: duty=105; 15'd15707: duty=115; 15'd15708: duty=89; 15'd15709: duty=85; 15'd15710: duty=95; 15'd15711: duty=83;
15'd15712: duty=95; 15'd15713: duty=97; 15'd15714: duty=97; 15'd15715: duty=73; 15'd15716: duty=69; 15'd15717: duty=74; 15'd15718: duty=81; 15'd15719: duty=94;
15'd15720: duty=77; 15'd15721: duty=78; 15'd15722: duty=93; 15'd15723: duty=89; 15'd15724: duty=100; 15'd15725: duty=102; 15'd15726: duty=103; 15'd15727: duty=106;
15'd15728: duty=105; 15'd15729: duty=114; 15'd15730: duty=103; 15'd15731: duty=99; 15'd15732: duty=106; 15'd15733: duty=108; 15'd15734: duty=110; 15'd15735: duty=114;
15'd15736: duty=118; 15'd15737: duty=135; 15'd15738: duty=124; 15'd15739: duty=116; 15'd15740: duty=133; 15'd15741: duty=128; 15'd15742: duty=134; 15'd15743: duty=146;
15'd15744: duty=147; 15'd15745: duty=140; 15'd15746: duty=148; 15'd15747: duty=151; 15'd15748: duty=151; 15'd15749: duty=157; 15'd15750: duty=170; 15'd15751: duty=178;
15'd15752: duty=175; 15'd15753: duty=181; 15'd15754: duty=174; 15'd15755: duty=170; 15'd15756: duty=164; 15'd15757: duty=162; 15'd15758: duty=160; 15'd15759: duty=169;
15'd15760: duty=182; 15'd15761: duty=177; 15'd15762: duty=170; 15'd15763: duty=179; 15'd15764: duty=179; 15'd15765: duty=173; 15'd15766: duty=185; 15'd15767: duty=180;
15'd15768: duty=178; 15'd15769: duty=190; 15'd15770: duty=188; 15'd15771: duty=185; 15'd15772: duty=176; 15'd15773: duty=168; 15'd15774: duty=157; 15'd15775: duty=148;
15'd15776: duty=146; 15'd15777: duty=144; 15'd15778: duty=145; 15'd15779: duty=128; 15'd15780: duty=127; 15'd15781: duty=127; 15'd15782: duty=120; 15'd15783: duty=113;
15'd15784: duty=98; 15'd15785: duty=94; 15'd15786: duty=98; 15'd15787: duty=107; 15'd15788: duty=110; 15'd15789: duty=108; 15'd15790: duty=98; 15'd15791: duty=93;
15'd15792: duty=92; 15'd15793: duty=82; 15'd15794: duty=90; 15'd15795: duty=107; 15'd15796: duty=87; 15'd15797: duty=78; 15'd15798: duty=80; 15'd15799: duty=82;
15'd15800: duty=90; 15'd15801: duty=92; 15'd15802: duty=81; 15'd15803: duty=73; 15'd15804: duty=102; 15'd15805: duty=93; 15'd15806: duty=83; 15'd15807: duty=90;
15'd15808: duty=88; 15'd15809: duty=87; 15'd15810: duty=81; 15'd15811: duty=83; 15'd15812: duty=93; 15'd15813: duty=109; 15'd15814: duty=110; 15'd15815: duty=106;
15'd15816: duty=111; 15'd15817: duty=114; 15'd15818: duty=111; 15'd15819: duty=112; 15'd15820: duty=120; 15'd15821: duty=135; 15'd15822: duty=145; 15'd15823: duty=142;
15'd15824: duty=125; 15'd15825: duty=127; 15'd15826: duty=135; 15'd15827: duty=135; 15'd15828: duty=145; 15'd15829: duty=153; 15'd15830: duty=169; 15'd15831: duty=155;
15'd15832: duty=155; 15'd15833: duty=153; 15'd15834: duty=154; 15'd15835: duty=176; 15'd15836: duty=163; 15'd15837: duty=173; 15'd15838: duty=181; 15'd15839: duty=184;
15'd15840: duty=203; 15'd15841: duty=197; 15'd15842: duty=180; 15'd15843: duty=173; 15'd15844: duty=171; 15'd15845: duty=178; 15'd15846: duty=175; 15'd15847: duty=173;
15'd15848: duty=183; 15'd15849: duty=170; 15'd15850: duty=164; 15'd15851: duty=164; 15'd15852: duty=166; 15'd15853: duty=184; 15'd15854: duty=166; 15'd15855: duty=157;
15'd15856: duty=155; 15'd15857: duty=149; 15'd15858: duty=155; 15'd15859: duty=158; 15'd15860: duty=154; 15'd15861: duty=145; 15'd15862: duty=148; 15'd15863: duty=124;
15'd15864: duty=118; 15'd15865: duty=125; 15'd15866: duty=127; 15'd15867: duty=113; 15'd15868: duty=107; 15'd15869: duty=113; 15'd15870: duty=110; 15'd15871: duty=111;
15'd15872: duty=103; 15'd15873: duty=80; 15'd15874: duty=75; 15'd15875: duty=86; 15'd15876: duty=86; 15'd15877: duty=94; 15'd15878: duty=94; 15'd15879: duty=91;
15'd15880: duty=86; 15'd15881: duty=88; 15'd15882: duty=93; 15'd15883: duty=97; 15'd15884: duty=88; 15'd15885: duty=90; 15'd15886: duty=93; 15'd15887: duty=90;
15'd15888: duty=76; 15'd15889: duty=84; 15'd15890: duty=97; 15'd15891: duty=84; 15'd15892: duty=82; 15'd15893: duty=96; 15'd15894: duty=118; 15'd15895: duty=127;
15'd15896: duty=116; 15'd15897: duty=103; 15'd15898: duty=99; 15'd15899: duty=108; 15'd15900: duty=114; 15'd15901: duty=116; 15'd15902: duty=118; 15'd15903: duty=112;
15'd15904: duty=120; 15'd15905: duty=120; 15'd15906: duty=140; 15'd15907: duty=141; 15'd15908: duty=138; 15'd15909: duty=138; 15'd15910: duty=136; 15'd15911: duty=143;
15'd15912: duty=138; 15'd15913: duty=136; 15'd15914: duty=140; 15'd15915: duty=152; 15'd15916: duty=149; 15'd15917: duty=149; 15'd15918: duty=155; 15'd15919: duty=152;
15'd15920: duty=161; 15'd15921: duty=162; 15'd15922: duty=164; 15'd15923: duty=166; 15'd15924: duty=182; 15'd15925: duty=174; 15'd15926: duty=172; 15'd15927: duty=175;
15'd15928: duty=166; 15'd15929: duty=175; 15'd15930: duty=191; 15'd15931: duty=191; 15'd15932: duty=189; 15'd15933: duty=190; 15'd15934: duty=186; 15'd15935: duty=195;
15'd15936: duty=197; 15'd15937: duty=183; 15'd15938: duty=160; 15'd15939: duty=161; 15'd15940: duty=154; 15'd15941: duty=154; 15'd15942: duty=145; 15'd15943: duty=136;
15'd15944: duty=138; 15'd15945: duty=147; 15'd15946: duty=142; 15'd15947: duty=134; 15'd15948: duty=124; 15'd15949: duty=134; 15'd15950: duty=137; 15'd15951: duty=137;
15'd15952: duty=139; 15'd15953: duty=136; 15'd15954: duty=123; 15'd15955: duty=114; 15'd15956: duty=98; 15'd15957: duty=107; 15'd15958: duty=120; 15'd15959: duty=107;
15'd15960: duty=99; 15'd15961: duty=91; 15'd15962: duty=92; 15'd15963: duty=83; 15'd15964: duty=96; 15'd15965: duty=74; 15'd15966: duty=67; 15'd15967: duty=84;
15'd15968: duty=81; 15'd15969: duty=74; 15'd15970: duty=84; 15'd15971: duty=84; 15'd15972: duty=83; 15'd15973: duty=82; 15'd15974: duty=86; 15'd15975: duty=86;
15'd15976: duty=110; 15'd15977: duty=101; 15'd15978: duty=101; 15'd15979: duty=99; 15'd15980: duty=87; 15'd15981: duty=96; 15'd15982: duty=104; 15'd15983: duty=104;
15'd15984: duty=101; 15'd15985: duty=106; 15'd15986: duty=96; 15'd15987: duty=101; 15'd15988: duty=121; 15'd15989: duty=129; 15'd15990: duty=129; 15'd15991: duty=125;
15'd15992: duty=128; 15'd15993: duty=139; 15'd15994: duty=123; 15'd15995: duty=131; 15'd15996: duty=137; 15'd15997: duty=143; 15'd15998: duty=141; 15'd15999: duty=151;
15'd16000: duty=146; 15'd16001: duty=160; 15'd16002: duty=159; 15'd16003: duty=162; 15'd16004: duty=158; 15'd16005: duty=166; 15'd16006: duty=173; 15'd16007: duty=158;
15'd16008: duty=159; 15'd16009: duty=161; 15'd16010: duty=158; 15'd16011: duty=178; 15'd16012: duty=184; 15'd16013: duty=168; 15'd16014: duty=188; 15'd16015: duty=186;
15'd16016: duty=185; 15'd16017: duty=198; 15'd16018: duty=191; 15'd16019: duty=178; 15'd16020: duty=189; 15'd16021: duty=171; 15'd16022: duty=157; 15'd16023: duty=155;
15'd16024: duty=170; 15'd16025: duty=161; 15'd16026: duty=149; 15'd16027: duty=146; 15'd16028: duty=146; 15'd16029: duty=144; 15'd16030: duty=135; 15'd16031: duty=132;
15'd16032: duty=131; 15'd16033: duty=135; 15'd16034: duty=127; 15'd16035: duty=125; 15'd16036: duty=133; 15'd16037: duty=131; 15'd16038: duty=119; 15'd16039: duty=108;
15'd16040: duty=100; 15'd16041: duty=109; 15'd16042: duty=112; 15'd16043: duty=102; 15'd16044: duty=98; 15'd16045: duty=96; 15'd16046: duty=104; 15'd16047: duty=97;
15'd16048: duty=95; 15'd16049: duty=104; 15'd16050: duty=93; 15'd16051: duty=98; 15'd16052: duty=101; 15'd16053: duty=82; 15'd16054: duty=92; 15'd16055: duty=94;
15'd16056: duty=78; 15'd16057: duty=96; 15'd16058: duty=91; 15'd16059: duty=95; 15'd16060: duty=99; 15'd16061: duty=97; 15'd16062: duty=98; 15'd16063: duty=111;
15'd16064: duty=124; 15'd16065: duty=112; 15'd16066: duty=115; 15'd16067: duty=118; 15'd16068: duty=121; 15'd16069: duty=124; 15'd16070: duty=125; 15'd16071: duty=124;
15'd16072: duty=107; 15'd16073: duty=121; 15'd16074: duty=112; 15'd16075: duty=102; 15'd16076: duty=122; 15'd16077: duty=124; 15'd16078: duty=127; 15'd16079: duty=131;
15'd16080: duty=136; 15'd16081: duty=139; 15'd16082: duty=145; 15'd16083: duty=146; 15'd16084: duty=159; 15'd16085: duty=151; 15'd16086: duty=154; 15'd16087: duty=170;
15'd16088: duty=169; 15'd16089: duty=163; 15'd16090: duty=164; 15'd16091: duty=170; 15'd16092: duty=171; 15'd16093: duty=168; 15'd16094: duty=156; 15'd16095: duty=165;
15'd16096: duty=177; 15'd16097: duty=177; 15'd16098: duty=166; 15'd16099: duty=170; 15'd16100: duty=183; 15'd16101: duty=180; 15'd16102: duty=179; 15'd16103: duty=170;
15'd16104: duty=170; 15'd16105: duty=176; 15'd16106: duty=159; 15'd16107: duty=154; 15'd16108: duty=156; 15'd16109: duty=151; 15'd16110: duty=150; 15'd16111: duty=131;
15'd16112: duty=141; 15'd16113: duty=143; 15'd16114: duty=133; 15'd16115: duty=133; 15'd16116: duty=124; 15'd16117: duty=131; 15'd16118: duty=124; 15'd16119: duty=122;
15'd16120: duty=112; 15'd16121: duty=90; 15'd16122: duty=110; 15'd16123: duty=108; 15'd16124: duty=101; 15'd16125: duty=106; 15'd16126: duty=87; 15'd16127: duty=92;
15'd16128: duty=89; 15'd16129: duty=105; 15'd16130: duty=112; 15'd16131: duty=102; 15'd16132: duty=96; 15'd16133: duty=85; 15'd16134: duty=90; 15'd16135: duty=102;
15'd16136: duty=88; 15'd16137: duty=85; 15'd16138: duty=87; 15'd16139: duty=84; 15'd16140: duty=98; 15'd16141: duty=87; 15'd16142: duty=89; 15'd16143: duty=96;
15'd16144: duty=93; 15'd16145: duty=87; 15'd16146: duty=99; 15'd16147: duty=125; 15'd16148: duty=122; 15'd16149: duty=110; 15'd16150: duty=101; 15'd16151: duty=102;
15'd16152: duty=104; 15'd16153: duty=104; 15'd16154: duty=104; 15'd16155: duty=105; 15'd16156: duty=139; 15'd16157: duty=143; 15'd16158: duty=138; 15'd16159: duty=142;
15'd16160: duty=150; 15'd16161: duty=148; 15'd16162: duty=131; 15'd16163: duty=139; 15'd16164: duty=158; 15'd16165: duty=152; 15'd16166: duty=147; 15'd16167: duty=145;
15'd16168: duty=139; 15'd16169: duty=157; 15'd16170: duty=157; 15'd16171: duty=169; 15'd16172: duty=174; 15'd16173: duty=183; 15'd16174: duty=185; 15'd16175: duty=180;
15'd16176: duty=184; 15'd16177: duty=188; 15'd16178: duty=181; 15'd16179: duty=171; 15'd16180: duty=174; 15'd16181: duty=179; 15'd16182: duty=187; 15'd16183: duty=176;
15'd16184: duty=175; 15'd16185: duty=189; 15'd16186: duty=188; 15'd16187: duty=179; 15'd16188: duty=183; 15'd16189: duty=185; 15'd16190: duty=182; 15'd16191: duty=166;
15'd16192: duty=150; 15'd16193: duty=151; 15'd16194: duty=143; 15'd16195: duty=137; 15'd16196: duty=142; 15'd16197: duty=121; 15'd16198: duty=116; 15'd16199: duty=124;
15'd16200: duty=117; 15'd16201: duty=109; 15'd16202: duty=104; 15'd16203: duty=107; 15'd16204: duty=102; 15'd16205: duty=100; 15'd16206: duty=96; 15'd16207: duty=95;
15'd16208: duty=90; 15'd16209: duty=80; 15'd16210: duty=73; 15'd16211: duty=85; 15'd16212: duty=90; 15'd16213: duty=81; 15'd16214: duty=82; 15'd16215: duty=87;
15'd16216: duty=85; 15'd16217: duty=71; 15'd16218: duty=76; 15'd16219: duty=93; 15'd16220: duty=93; 15'd16221: duty=90; 15'd16222: duty=91; 15'd16223: duty=102;
15'd16224: duty=89; 15'd16225: duty=84; 15'd16226: duty=97; 15'd16227: duty=100; 15'd16228: duty=95; 15'd16229: duty=91; 15'd16230: duty=121; 15'd16231: duty=108;
15'd16232: duty=112; 15'd16233: duty=113; 15'd16234: duty=115; 15'd16235: duty=132; 15'd16236: duty=128; 15'd16237: duty=125; 15'd16238: duty=118; 15'd16239: duty=119;
15'd16240: duty=131; 15'd16241: duty=140; 15'd16242: duty=130; 15'd16243: duty=134; 15'd16244: duty=155; 15'd16245: duty=157; 15'd16246: duty=158; 15'd16247: duty=154;
15'd16248: duty=141; 15'd16249: duty=148; 15'd16250: duty=148; 15'd16251: duty=155; 15'd16252: duty=153; 15'd16253: duty=146; 15'd16254: duty=144; 15'd16255: duty=151;
15'd16256: duty=147; 15'd16257: duty=153; 15'd16258: duty=171; 15'd16259: duty=176; 15'd16260: duty=168; 15'd16261: duty=160; 15'd16262: duty=171; 15'd16263: duty=179;
15'd16264: duty=186; 15'd16265: duty=190; 15'd16266: duty=185; 15'd16267: duty=176; 15'd16268: duty=181; 15'd16269: duty=184; 15'd16270: duty=184; 15'd16271: duty=185;
15'd16272: duty=170; 15'd16273: duty=156; 15'd16274: duty=159; 15'd16275: duty=157; 15'd16276: duty=157; 15'd16277: duty=157; 15'd16278: duty=140; 15'd16279: duty=143;
15'd16280: duty=135; 15'd16281: duty=143; 15'd16282: duty=137; 15'd16283: duty=121; 15'd16284: duty=120; 15'd16285: duty=116; 15'd16286: duty=124; 15'd16287: duty=111;
15'd16288: duty=115; 15'd16289: duty=111; 15'd16290: duty=104; 15'd16291: duty=97; 15'd16292: duty=100; 15'd16293: duty=100; 15'd16294: duty=91; 15'd16295: duty=97;
15'd16296: duty=94; 15'd16297: duty=77; 15'd16298: duty=82; 15'd16299: duty=81; 15'd16300: duty=74; 15'd16301: duty=78; 15'd16302: duty=88; 15'd16303: duty=104;
15'd16304: duty=94; 15'd16305: duty=81; 15'd16306: duty=82; 15'd16307: duty=92; 15'd16308: duty=98; 15'd16309: duty=106; 15'd16310: duty=97; 15'd16311: duty=103;
15'd16312: duty=111; 15'd16313: duty=106; 15'd16314: duty=115; 15'd16315: duty=115; 15'd16316: duty=117; 15'd16317: duty=129; 15'd16318: duty=119; 15'd16319: duty=114;
15'd16320: duty=114; 15'd16321: duty=114; 15'd16322: duty=120; 15'd16323: duty=106; 15'd16324: duty=111; 15'd16325: duty=128; 15'd16326: duty=140; 15'd16327: duty=156;
15'd16328: duty=155; 15'd16329: duty=144; 15'd16330: duty=165; 15'd16331: duty=157; 15'd16332: duty=153; 15'd16333: duty=163; 15'd16334: duty=155; 15'd16335: duty=152;
15'd16336: duty=135; 15'd16337: duty=136; 15'd16338: duty=155; 15'd16339: duty=163; 15'd16340: duty=164; 15'd16341: duty=169; 15'd16342: duty=170; 15'd16343: duty=174;
15'd16344: duty=172; 15'd16345: duty=180; 15'd16346: duty=172; 15'd16347: duty=180; 15'd16348: duty=187; 15'd16349: duty=180; 15'd16350: duty=187; 15'd16351: duty=191;
15'd16352: duty=190; 15'd16353: duty=174; 15'd16354: duty=165; 15'd16355: duty=164; 15'd16356: duty=169; 15'd16357: duty=146; 15'd16358: duty=146; 15'd16359: duty=141;
15'd16360: duty=144; 15'd16361: duty=141; 15'd16362: duty=118; 15'd16363: duty=126; 15'd16364: duty=132; 15'd16365: duty=123; 15'd16366: duty=114; 15'd16367: duty=117;
15'd16368: duty=125; 15'd16369: duty=126; 15'd16370: duty=112; 15'd16371: duty=107; 15'd16372: duty=101; 15'd16373: duty=99; 15'd16374: duty=103; 15'd16375: duty=96;
15'd16376: duty=92; 15'd16377: duty=93; 15'd16378: duty=90; 15'd16379: duty=82; 15'd16380: duty=75; 15'd16381: duty=84; 15'd16382: duty=96; 15'd16383: duty=84;
15'd16384: duty=84; 15'd16385: duty=94; 15'd16386: duty=92; 15'd16387: duty=90; 15'd16388: duty=81; 15'd16389: duty=96; 15'd16390: duty=99; 15'd16391: duty=93;
15'd16392: duty=84; 15'd16393: duty=84; 15'd16394: duty=107; 15'd16395: duty=112; 15'd16396: duty=116; 15'd16397: duty=109; 15'd16398: duty=107; 15'd16399: duty=124;
15'd16400: duty=134; 15'd16401: duty=141; 15'd16402: duty=125; 15'd16403: duty=123; 15'd16404: duty=125; 15'd16405: duty=121; 15'd16406: duty=127; 15'd16407: duty=121;
15'd16408: duty=137; 15'd16409: duty=144; 15'd16410: duty=139; 15'd16411: duty=141; 15'd16412: duty=136; 15'd16413: duty=140; 15'd16414: duty=149; 15'd16415: duty=153;
15'd16416: duty=154; 15'd16417: duty=160; 15'd16418: duty=162; 15'd16419: duty=165; 15'd16420: duty=157; 15'd16421: duty=163; 15'd16422: duty=166; 15'd16423: duty=158;
15'd16424: duty=166; 15'd16425: duty=171; 15'd16426: duty=188; 15'd16427: duty=176; 15'd16428: duty=191; 15'd16429: duty=196; 15'd16430: duty=184; 15'd16431: duty=177;
15'd16432: duty=182; 15'd16433: duty=180; 15'd16434: duty=168; 15'd16435: duty=166; 15'd16436: duty=165; 15'd16437: duty=167; 15'd16438: duty=157; 15'd16439: duty=150;
15'd16440: duty=142; 15'd16441: duty=145; 15'd16442: duty=142; 15'd16443: duty=145; 15'd16444: duty=139; 15'd16445: duty=131; 15'd16446: duty=127; 15'd16447: duty=139;
15'd16448: duty=146; 15'd16449: duty=133; 15'd16450: duty=113; 15'd16451: duty=99; 15'd16452: duty=108; 15'd16453: duty=121; 15'd16454: duty=120; 15'd16455: duty=123;
15'd16456: duty=107; 15'd16457: duty=100; 15'd16458: duty=90; 15'd16459: duty=86; 15'd16460: duty=96; 15'd16461: duty=90; 15'd16462: duty=88; 15'd16463: duty=87;
15'd16464: duty=76; 15'd16465: duty=86; 15'd16466: duty=96; 15'd16467: duty=98; 15'd16468: duty=87; 15'd16469: duty=95; 15'd16470: duty=108; 15'd16471: duty=101;
15'd16472: duty=113; 15'd16473: duty=101; 15'd16474: duty=88; 15'd16475: duty=84; 15'd16476: duty=81; 15'd16477: duty=84; 15'd16478: duty=109; 15'd16479: duty=109;
15'd16480: duty=112; 15'd16481: duty=107; 15'd16482: duty=108; 15'd16483: duty=110; 15'd16484: duty=121; 15'd16485: duty=124; 15'd16486: duty=107; 15'd16487: duty=119;
15'd16488: duty=128; 15'd16489: duty=131; 15'd16490: duty=140; 15'd16491: duty=137; 15'd16492: duty=138; 15'd16493: duty=153; 15'd16494: duty=145; 15'd16495: duty=142;
15'd16496: duty=151; 15'd16497: duty=151; 15'd16498: duty=163; 15'd16499: duty=163; 15'd16500: duty=148; 15'd16501: duty=155; 15'd16502: duty=159; 15'd16503: duty=163;
15'd16504: duty=165; 15'd16505: duty=162; 15'd16506: duty=164; 15'd16507: duty=171; 15'd16508: duty=168; 15'd16509: duty=163; 15'd16510: duty=167; 15'd16511: duty=180;
15'd16512: duty=176; 15'd16513: duty=165; 15'd16514: duty=175; 15'd16515: duty=181; 15'd16516: duty=180; 15'd16517: duty=173; 15'd16518: duty=165; 15'd16519: duty=172;
15'd16520: duty=167; 15'd16521: duty=160; 15'd16522: duty=155; 15'd16523: duty=146; 15'd16524: duty=146; 15'd16525: duty=145; 15'd16526: duty=144; 15'd16527: duty=146;
15'd16528: duty=147; 15'd16529: duty=139; 15'd16530: duty=127; 15'd16531: duty=136; 15'd16532: duty=131; 15'd16533: duty=121; 15'd16534: duty=119; 15'd16535: duty=103;
15'd16536: duty=110; 15'd16537: duty=116; 15'd16538: duty=110; 15'd16539: duty=98; 15'd16540: duty=95; 15'd16541: duty=96; 15'd16542: duty=94; 15'd16543: duty=90;
15'd16544: duty=95; 15'd16545: duty=92; 15'd16546: duty=91; 15'd16547: duty=105; 15'd16548: duty=88; 15'd16549: duty=79; 15'd16550: duty=90; 15'd16551: duty=93;
15'd16552: duty=94; 15'd16553: duty=99; 15'd16554: duty=102; 15'd16555: duty=98; 15'd16556: duty=101; 15'd16557: duty=106; 15'd16558: duty=94; 15'd16559: duty=95;
15'd16560: duty=111; 15'd16561: duty=104; 15'd16562: duty=108; 15'd16563: duty=113; 15'd16564: duty=119; 15'd16565: duty=137; 15'd16566: duty=111; 15'd16567: duty=110;
15'd16568: duty=111; 15'd16569: duty=106; 15'd16570: duty=121; 15'd16571: duty=124; 15'd16572: duty=127; 15'd16573: duty=124; 15'd16574: duty=119; 15'd16575: duty=115;
15'd16576: duty=131; 15'd16577: duty=152; 15'd16578: duty=151; 15'd16579: duty=144; 15'd16580: duty=149; 15'd16581: duty=144; 15'd16582: duty=151; 15'd16583: duty=160;
15'd16584: duty=140; 15'd16585: duty=153; 15'd16586: duty=162; 15'd16587: duty=157; 15'd16588: duty=160; 15'd16589: duty=156; 15'd16590: duty=157; 15'd16591: duty=151;
15'd16592: duty=152; 15'd16593: duty=157; 15'd16594: duty=168; 15'd16595: duty=173; 15'd16596: duty=177; 15'd16597: duty=182; 15'd16598: duty=188; 15'd16599: duty=185;
15'd16600: duty=190; 15'd16601: duty=189; 15'd16602: duty=185; 15'd16603: duty=186; 15'd16604: duty=177; 15'd16605: duty=169; 15'd16606: duty=161; 15'd16607: duty=160;
15'd16608: duty=155; 15'd16609: duty=152; 15'd16610: duty=147; 15'd16611: duty=147; 15'd16612: duty=143; 15'd16613: duty=138; 15'd16614: duty=130; 15'd16615: duty=134;
15'd16616: duty=135; 15'd16617: duty=133; 15'd16618: duty=129; 15'd16619: duty=117; 15'd16620: duty=111; 15'd16621: duty=112; 15'd16622: duty=104; 15'd16623: duty=94;
15'd16624: duty=89; 15'd16625: duty=94; 15'd16626: duty=102; 15'd16627: duty=106; 15'd16628: duty=100; 15'd16629: duty=103; 15'd16630: duty=88; 15'd16631: duty=81;
15'd16632: duty=87; 15'd16633: duty=86; 15'd16634: duty=99; 15'd16635: duty=81; 15'd16636: duty=73; 15'd16637: duty=70; 15'd16638: duty=73; 15'd16639: duty=78;
15'd16640: duty=91; 15'd16641: duty=90; 15'd16642: duty=87; 15'd16643: duty=93; 15'd16644: duty=95; 15'd16645: duty=93; 15'd16646: duty=97; 15'd16647: duty=104;
15'd16648: duty=97; 15'd16649: duty=102; 15'd16650: duty=114; 15'd16651: duty=113; 15'd16652: duty=107; 15'd16653: duty=98; 15'd16654: duty=119; 15'd16655: duty=128;
15'd16656: duty=132; 15'd16657: duty=137; 15'd16658: duty=138; 15'd16659: duty=151; 15'd16660: duty=144; 15'd16661: duty=141; 15'd16662: duty=142; 15'd16663: duty=146;
15'd16664: duty=152; 15'd16665: duty=148; 15'd16666: duty=146; 15'd16667: duty=142; 15'd16668: duty=155; 15'd16669: duty=171; 15'd16670: duty=162; 15'd16671: duty=169;
15'd16672: duty=170; 15'd16673: duty=177; 15'd16674: duty=185; 15'd16675: duty=196; 15'd16676: duty=192; 15'd16677: duty=186; 15'd16678: duty=179; 15'd16679: duty=175;
15'd16680: duty=179; 15'd16681: duty=185; 15'd16682: duty=186; 15'd16683: duty=182; 15'd16684: duty=180; 15'd16685: duty=185; 15'd16686: duty=180; 15'd16687: duty=174;
15'd16688: duty=169; 15'd16689: duty=174; 15'd16690: duty=160; 15'd16691: duty=162; 15'd16692: duty=163; 15'd16693: duty=153; 15'd16694: duty=153; 15'd16695: duty=147;
15'd16696: duty=147; 15'd16697: duty=133; 15'd16698: duty=130; 15'd16699: duty=125; 15'd16700: duty=124; 15'd16701: duty=117; 15'd16702: duty=119; 15'd16703: duty=112;
15'd16704: duty=100; 15'd16705: duty=84; 15'd16706: duty=86; 15'd16707: duty=81; 15'd16708: duty=90; 15'd16709: duty=95; 15'd16710: duty=90; 15'd16711: duty=81;
15'd16712: duty=91; 15'd16713: duty=82; 15'd16714: duty=76; 15'd16715: duty=82; 15'd16716: duty=89; 15'd16717: duty=84; 15'd16718: duty=77; 15'd16719: duty=79;
15'd16720: duty=64; 15'd16721: duty=84; 15'd16722: duty=84; 15'd16723: duty=74; 15'd16724: duty=89; 15'd16725: duty=96; 15'd16726: duty=86; 15'd16727: duty=98;
15'd16728: duty=101; 15'd16729: duty=99; 15'd16730: duty=98; 15'd16731: duty=114; 15'd16732: duty=113; 15'd16733: duty=121; 15'd16734: duty=127; 15'd16735: duty=128;
15'd16736: duty=130; 15'd16737: duty=135; 15'd16738: duty=131; 15'd16739: duty=133; 15'd16740: duty=151; 15'd16741: duty=131; 15'd16742: duty=133; 15'd16743: duty=137;
15'd16744: duty=124; 15'd16745: duty=139; 15'd16746: duty=150; 15'd16747: duty=143; 15'd16748: duty=150; 15'd16749: duty=152; 15'd16750: duty=158; 15'd16751: duty=151;
15'd16752: duty=159; 15'd16753: duty=173; 15'd16754: duty=168; 15'd16755: duty=185; 15'd16756: duty=193; 15'd16757: duty=185; 15'd16758: duty=186; 15'd16759: duty=184;
15'd16760: duty=174; 15'd16761: duty=179; 15'd16762: duty=182; 15'd16763: duty=181; 15'd16764: duty=177; 15'd16765: duty=175; 15'd16766: duty=169; 15'd16767: duty=168;
15'd16768: duty=167; 15'd16769: duty=155; 15'd16770: duty=151; 15'd16771: duty=145; 15'd16772: duty=146; 15'd16773: duty=145; 15'd16774: duty=141; 15'd16775: duty=130;
15'd16776: duty=141; 15'd16777: duty=150; 15'd16778: duty=144; 15'd16779: duty=141; 15'd16780: duty=146; 15'd16781: duty=130; 15'd16782: duty=128; 15'd16783: duty=117;
15'd16784: duty=112; 15'd16785: duty=107; 15'd16786: duty=105; 15'd16787: duty=103; 15'd16788: duty=102; 15'd16789: duty=106; 15'd16790: duty=98; 15'd16791: duty=93;
15'd16792: duty=97; 15'd16793: duty=103; 15'd16794: duty=93; 15'd16795: duty=102; 15'd16796: duty=108; 15'd16797: duty=102; 15'd16798: duty=96; 15'd16799: duty=108;
15'd16800: duty=93; 15'd16801: duty=99; 15'd16802: duty=102; 15'd16803: duty=101; 15'd16804: duty=99; 15'd16805: duty=107; 15'd16806: duty=108; 15'd16807: duty=105;
15'd16808: duty=104; 15'd16809: duty=99; 15'd16810: duty=98; 15'd16811: duty=102; 15'd16812: duty=113; 15'd16813: duty=114; 15'd16814: duty=119; 15'd16815: duty=111;
15'd16816: duty=117; 15'd16817: duty=129; 15'd16818: duty=120; 15'd16819: duty=109; 15'd16820: duty=121; 15'd16821: duty=134; 15'd16822: duty=126; 15'd16823: duty=131;
15'd16824: duty=141; 15'd16825: duty=125; 15'd16826: duty=119; 15'd16827: duty=119; 15'd16828: duty=118; 15'd16829: duty=133; 15'd16830: duty=145; 15'd16831: duty=143;
15'd16832: duty=143; 15'd16833: duty=139; 15'd16834: duty=146; 15'd16835: duty=154; 15'd16836: duty=152; 15'd16837: duty=153; 15'd16838: duty=163; 15'd16839: duty=164;
15'd16840: duty=163; 15'd16841: duty=164; 15'd16842: duty=169; 15'd16843: duty=167; 15'd16844: duty=172; 15'd16845: duty=176; 15'd16846: duty=163; 15'd16847: duty=162;
15'd16848: duty=172; 15'd16849: duty=176; 15'd16850: duty=178; 15'd16851: duty=176; 15'd16852: duty=176; 15'd16853: duty=173; 15'd16854: duty=157; 15'd16855: duty=158;
15'd16856: duty=153; 15'd16857: duty=144; 15'd16858: duty=143; 15'd16859: duty=144; 15'd16860: duty=148; 15'd16861: duty=140; 15'd16862: duty=132; 15'd16863: duty=140;
15'd16864: duty=130; 15'd16865: duty=133; 15'd16866: duty=137; 15'd16867: duty=137; 15'd16868: duty=122; 15'd16869: duty=119; 15'd16870: duty=124; 15'd16871: duty=113;
15'd16872: duty=102; 15'd16873: duty=96; 15'd16874: duty=105; 15'd16875: duty=107; 15'd16876: duty=107; 15'd16877: duty=97; 15'd16878: duty=95; 15'd16879: duty=102;
15'd16880: duty=99; 15'd16881: duty=91; 15'd16882: duty=95; 15'd16883: duty=106; 15'd16884: duty=112; 15'd16885: duty=110; 15'd16886: duty=110; 15'd16887: duty=104;
15'd16888: duty=106; 15'd16889: duty=122; 15'd16890: duty=110; 15'd16891: duty=94; 15'd16892: duty=94; 15'd16893: duty=96; 15'd16894: duty=105; 15'd16895: duty=106;
15'd16896: duty=105; 15'd16897: duty=121; 15'd16898: duty=121; 15'd16899: duty=106; 15'd16900: duty=104; 15'd16901: duty=110; 15'd16902: duty=111; 15'd16903: duty=119;
15'd16904: duty=125; 15'd16905: duty=121; 15'd16906: duty=124; 15'd16907: duty=143; 15'd16908: duty=144; 15'd16909: duty=124; 15'd16910: duty=121; 15'd16911: duty=130;
15'd16912: duty=132; 15'd16913: duty=133; 15'd16914: duty=134; 15'd16915: duty=135; 15'd16916: duty=135; 15'd16917: duty=129; 15'd16918: duty=127; 15'd16919: duty=130;
15'd16920: duty=146; 15'd16921: duty=150; 15'd16922: duty=155; 15'd16923: duty=165; 15'd16924: duty=163; 15'd16925: duty=161; 15'd16926: duty=155; 15'd16927: duty=162;
15'd16928: duty=172; 15'd16929: duty=185; 15'd16930: duty=185; 15'd16931: duty=180; 15'd16932: duty=179; 15'd16933: duty=176; 15'd16934: duty=182; 15'd16935: duty=173;
15'd16936: duty=159; 15'd16937: duty=172; 15'd16938: duty=167; 15'd16939: duty=152; 15'd16940: duty=147; 15'd16941: duty=141; 15'd16942: duty=145; 15'd16943: duty=148;
15'd16944: duty=140; 15'd16945: duty=142; 15'd16946: duty=142; 15'd16947: duty=145; 15'd16948: duty=148; 15'd16949: duty=139; 15'd16950: duty=131; 15'd16951: duty=118;
15'd16952: duty=113; 15'd16953: duty=107; 15'd16954: duty=104; 15'd16955: duty=116; 15'd16956: duty=105; 15'd16957: duty=108; 15'd16958: duty=116; 15'd16959: duty=109;
15'd16960: duty=107; 15'd16961: duty=97; 15'd16962: duty=96; 15'd16963: duty=99; 15'd16964: duty=99; 15'd16965: duty=94; 15'd16966: duty=101; 15'd16967: duty=107;
15'd16968: duty=108; 15'd16969: duty=106; 15'd16970: duty=97; 15'd16971: duty=86; 15'd16972: duty=91; 15'd16973: duty=93; 15'd16974: duty=105; 15'd16975: duty=106;
15'd16976: duty=102; 15'd16977: duty=101; 15'd16978: duty=112; 15'd16979: duty=123; 15'd16980: duty=92; 15'd16981: duty=108; 15'd16982: duty=118; 15'd16983: duty=119;
15'd16984: duty=116; 15'd16985: duty=101; 15'd16986: duty=109; 15'd16987: duty=119; 15'd16988: duty=118; 15'd16989: duty=128; 15'd16990: duty=133; 15'd16991: duty=135;
15'd16992: duty=146; 15'd16993: duty=137; 15'd16994: duty=149; 15'd16995: duty=140; 15'd16996: duty=125; 15'd16997: duty=138; 15'd16998: duty=141; 15'd16999: duty=147;
15'd17000: duty=144; 15'd17001: duty=137; 15'd17002: duty=139; 15'd17003: duty=143; 15'd17004: duty=158; 15'd17005: duty=166; 15'd17006: duty=172; 15'd17007: duty=173;
15'd17008: duty=164; 15'd17009: duty=173; 15'd17010: duty=177; 15'd17011: duty=166; 15'd17012: duty=167; 15'd17013: duty=169; 15'd17014: duty=174; 15'd17015: duty=182;
15'd17016: duty=187; 15'd17017: duty=179; 15'd17018: duty=174; 15'd17019: duty=172; 15'd17020: duty=164; 15'd17021: duty=157; 15'd17022: duty=155; 15'd17023: duty=153;
15'd17024: duty=144; 15'd17025: duty=151; 15'd17026: duty=144; 15'd17027: duty=139; 15'd17028: duty=144; 15'd17029: duty=137; 15'd17030: duty=142; 15'd17031: duty=133;
15'd17032: duty=130; 15'd17033: duty=134; 15'd17034: duty=127; 15'd17035: duty=119; 15'd17036: duty=106; 15'd17037: duty=105; 15'd17038: duty=107; 15'd17039: duty=98;
15'd17040: duty=104; 15'd17041: duty=102; 15'd17042: duty=95; 15'd17043: duty=94; 15'd17044: duty=98; 15'd17045: duty=98; 15'd17046: duty=82; 15'd17047: duty=94;
15'd17048: duty=104; 15'd17049: duty=101; 15'd17050: duty=95; 15'd17051: duty=92; 15'd17052: duty=92; 15'd17053: duty=90; 15'd17054: duty=82; 15'd17055: duty=84;
15'd17056: duty=84; 15'd17057: duty=98; 15'd17058: duty=99; 15'd17059: duty=91; 15'd17060: duty=103; 15'd17061: duty=93; 15'd17062: duty=107; 15'd17063: duty=120;
15'd17064: duty=128; 15'd17065: duty=125; 15'd17066: duty=124; 15'd17067: duty=122; 15'd17068: duty=120; 15'd17069: duty=117; 15'd17070: duty=117; 15'd17071: duty=124;
15'd17072: duty=114; 15'd17073: duty=110; 15'd17074: duty=118; 15'd17075: duty=126; 15'd17076: duty=142; 15'd17077: duty=134; 15'd17078: duty=137; 15'd17079: duty=153;
15'd17080: duty=153; 15'd17081: duty=154; 15'd17082: duty=151; 15'd17083: duty=167; 15'd17084: duty=152; 15'd17085: duty=152; 15'd17086: duty=165; 15'd17087: duty=164;
15'd17088: duty=170; 15'd17089: duty=178; 15'd17090: duty=171; 15'd17091: duty=168; 15'd17092: duty=173; 15'd17093: duty=180; 15'd17094: duty=174; 15'd17095: duty=166;
15'd17096: duty=178; 15'd17097: duty=182; 15'd17098: duty=189; 15'd17099: duty=185; 15'd17100: duty=170; 15'd17101: duty=161; 15'd17102: duty=163; 15'd17103: duty=160;
15'd17104: duty=162; 15'd17105: duty=159; 15'd17106: duty=143; 15'd17107: duty=138; 15'd17108: duty=136; 15'd17109: duty=132; 15'd17110: duty=131; 15'd17111: duty=140;
15'd17112: duty=140; 15'd17113: duty=133; 15'd17114: duty=128; 15'd17115: duty=124; 15'd17116: duty=122; 15'd17117: duty=115; 15'd17118: duty=119; 15'd17119: duty=113;
15'd17120: duty=116; 15'd17121: duty=118; 15'd17122: duty=112; 15'd17123: duty=104; 15'd17124: duty=91; 15'd17125: duty=87; 15'd17126: duty=90; 15'd17127: duty=92;
15'd17128: duty=87; 15'd17129: duty=95; 15'd17130: duty=96; 15'd17131: duty=96; 15'd17132: duty=94; 15'd17133: duty=80; 15'd17134: duty=102; 15'd17135: duty=104;
15'd17136: duty=94; 15'd17137: duty=104; 15'd17138: duty=96; 15'd17139: duty=103; 15'd17140: duty=107; 15'd17141: duty=104; 15'd17142: duty=95; 15'd17143: duty=93;
15'd17144: duty=100; 15'd17145: duty=104; 15'd17146: duty=118; 15'd17147: duty=123; 15'd17148: duty=119; 15'd17149: duty=118; 15'd17150: duty=119; 15'd17151: duty=114;
15'd17152: duty=125; 15'd17153: duty=127; 15'd17154: duty=124; 15'd17155: duty=140; 15'd17156: duty=137; 15'd17157: duty=139; 15'd17158: duty=136; 15'd17159: duty=136;
15'd17160: duty=131; 15'd17161: duty=144; 15'd17162: duty=160; 15'd17163: duty=156; 15'd17164: duty=160; 15'd17165: duty=157; 15'd17166: duty=145; 15'd17167: duty=142;
15'd17168: duty=157; 15'd17169: duty=167; 15'd17170: duty=169; 15'd17171: duty=165; 15'd17172: duty=154; 15'd17173: duty=170; 15'd17174: duty=171; 15'd17175: duty=174;
15'd17176: duty=175; 15'd17177: duty=169; 15'd17178: duty=177; 15'd17179: duty=170; 15'd17180: duty=162; 15'd17181: duty=168; 15'd17182: duty=172; 15'd17183: duty=166;
15'd17184: duty=166; 15'd17185: duty=168; 15'd17186: duty=165; 15'd17187: duty=152; 15'd17188: duty=149; 15'd17189: duty=138; 15'd17190: duty=140; 15'd17191: duty=135;
15'd17192: duty=131; 15'd17193: duty=132; 15'd17194: duty=119; 15'd17195: duty=123; 15'd17196: duty=129; 15'd17197: duty=120; 15'd17198: duty=120; 15'd17199: duty=125;
15'd17200: duty=117; 15'd17201: duty=109; 15'd17202: duty=98; 15'd17203: duty=96; 15'd17204: duty=100; 15'd17205: duty=96; 15'd17206: duty=98; 15'd17207: duty=97;
15'd17208: duty=81; 15'd17209: duty=83; 15'd17210: duty=81; 15'd17211: duty=96; 15'd17212: duty=92; 15'd17213: duty=85; 15'd17214: duty=92; 15'd17215: duty=96;
15'd17216: duty=97; 15'd17217: duty=96; 15'd17218: duty=112; 15'd17219: duty=101; 15'd17220: duty=92; 15'd17221: duty=98; 15'd17222: duty=102; 15'd17223: duty=114;
15'd17224: duty=118; 15'd17225: duty=115; 15'd17226: duty=109; 15'd17227: duty=115; 15'd17228: duty=134; 15'd17229: duty=136; 15'd17230: duty=117; 15'd17231: duty=118;
15'd17232: duty=125; 15'd17233: duty=124; 15'd17234: duty=136; 15'd17235: duty=131; 15'd17236: duty=140; 15'd17237: duty=141; 15'd17238: duty=135; 15'd17239: duty=144;
15'd17240: duty=149; 15'd17241: duty=149; 15'd17242: duty=149; 15'd17243: duty=145; 15'd17244: duty=157; 15'd17245: duty=155; 15'd17246: duty=157; 15'd17247: duty=158;
15'd17248: duty=139; 15'd17249: duty=151; 15'd17250: duty=156; 15'd17251: duty=151; 15'd17252: duty=160; 15'd17253: duty=159; 15'd17254: duty=158; 15'd17255: duty=174;
15'd17256: duty=171; 15'd17257: duty=172; 15'd17258: duty=170; 15'd17259: duty=171; 15'd17260: duty=175; 15'd17261: duty=177; 15'd17262: duty=180; 15'd17263: duty=179;
15'd17264: duty=167; 15'd17265: duty=159; 15'd17266: duty=160; 15'd17267: duty=157; 15'd17268: duty=142; 15'd17269: duty=147; 15'd17270: duty=146; 15'd17271: duty=138;
15'd17272: duty=137; 15'd17273: duty=136; 15'd17274: duty=135; 15'd17275: duty=130; 15'd17276: duty=138; 15'd17277: duty=144; 15'd17278: duty=142; 15'd17279: duty=128;
15'd17280: duty=128; 15'd17281: duty=116; 15'd17282: duty=107; 15'd17283: duty=101; 15'd17284: duty=98; 15'd17285: duty=100; 15'd17286: duty=108; 15'd17287: duty=92;
15'd17288: duty=90; 15'd17289: duty=102; 15'd17290: duty=101; 15'd17291: duty=93; 15'd17292: duty=87; 15'd17293: duty=86; 15'd17294: duty=88; 15'd17295: duty=95;
15'd17296: duty=104; 15'd17297: duty=108; 15'd17298: duty=84; 15'd17299: duty=76; 15'd17300: duty=98; 15'd17301: duty=102; 15'd17302: duty=99; 15'd17303: duty=96;
15'd17304: duty=93; 15'd17305: duty=96; 15'd17306: duty=84; 15'd17307: duty=89; 15'd17308: duty=97; 15'd17309: duty=111; 15'd17310: duty=110; 15'd17311: duty=114;
15'd17312: duty=130; 15'd17313: duty=125; 15'd17314: duty=127; 15'd17315: duty=132; 15'd17316: duty=112; 15'd17317: duty=128; 15'd17318: duty=143; 15'd17319: duty=141;
15'd17320: duty=146; 15'd17321: duty=140; 15'd17322: duty=132; 15'd17323: duty=122; 15'd17324: duty=129; 15'd17325: duty=150; 15'd17326: duty=144; 15'd17327: duty=146;
15'd17328: duty=145; 15'd17329: duty=149; 15'd17330: duty=152; 15'd17331: duty=144; 15'd17332: duty=155; 15'd17333: duty=169; 15'd17334: duty=162; 15'd17335: duty=157;
15'd17336: duty=169; 15'd17337: duty=168; 15'd17338: duty=183; 15'd17339: duty=177; 15'd17340: duty=172; 15'd17341: duty=165; 15'd17342: duty=166; 15'd17343: duty=182;
15'd17344: duty=188; 15'd17345: duty=174; 15'd17346: duty=182; 15'd17347: duty=177; 15'd17348: duty=174; 15'd17349: duty=182; 15'd17350: duty=175; 15'd17351: duty=167;
15'd17352: duty=152; 15'd17353: duty=158; 15'd17354: duty=162; 15'd17355: duty=146; 15'd17356: duty=149; 15'd17357: duty=141; 15'd17358: duty=132; 15'd17359: duty=135;
15'd17360: duty=130; 15'd17361: duty=127; 15'd17362: duty=120; 15'd17363: duty=112; 15'd17364: duty=114; 15'd17365: duty=109; 15'd17366: duty=105; 15'd17367: duty=106;
15'd17368: duty=103; 15'd17369: duty=107; 15'd17370: duty=97; 15'd17371: duty=101; 15'd17372: duty=102; 15'd17373: duty=95; 15'd17374: duty=93; 15'd17375: duty=87;
15'd17376: duty=85; 15'd17377: duty=102; 15'd17378: duty=92; 15'd17379: duty=98; 15'd17380: duty=98; 15'd17381: duty=85; 15'd17382: duty=86; 15'd17383: duty=108;
15'd17384: duty=112; 15'd17385: duty=107; 15'd17386: duty=102; 15'd17387: duty=90; 15'd17388: duty=95; 15'd17389: duty=94; 15'd17390: duty=117; 15'd17391: duty=108;
15'd17392: duty=99; 15'd17393: duty=108; 15'd17394: duty=100; 15'd17395: duty=105; 15'd17396: duty=122; 15'd17397: duty=115; 15'd17398: duty=110; 15'd17399: duty=117;
15'd17400: duty=120; 15'd17401: duty=120; 15'd17402: duty=138; 15'd17403: duty=135; 15'd17404: duty=127; 15'd17405: duty=132; 15'd17406: duty=129; 15'd17407: duty=131;
15'd17408: duty=144; 15'd17409: duty=152; 15'd17410: duty=142; 15'd17411: duty=127; 15'd17412: duty=130; 15'd17413: duty=135; 15'd17414: duty=147; 15'd17415: duty=160;
15'd17416: duty=148; 15'd17417: duty=155; 15'd17418: duty=167; 15'd17419: duty=172; 15'd17420: duty=174; 15'd17421: duty=182; 15'd17422: duty=179; 15'd17423: duty=163;
15'd17424: duty=176; 15'd17425: duty=180; 15'd17426: duty=174; 15'd17427: duty=187; 15'd17428: duty=184; 15'd17429: duty=174; 15'd17430: duty=180; 15'd17431: duty=173;
15'd17432: duty=170; 15'd17433: duty=165; 15'd17434: duty=154; 15'd17435: duty=152; 15'd17436: duty=153; 15'd17437: duty=149; 15'd17438: duty=139; 15'd17439: duty=136;
15'd17440: duty=141; 15'd17441: duty=145; 15'd17442: duty=139; 15'd17443: duty=137; 15'd17444: duty=139; 15'd17445: duty=143; 15'd17446: duty=141; 15'd17447: duty=132;
15'd17448: duty=128; 15'd17449: duty=121; 15'd17450: duty=116; 15'd17451: duty=107; 15'd17452: duty=99; 15'd17453: duty=110; 15'd17454: duty=107; 15'd17455: duty=98;
15'd17456: duty=81; 15'd17457: duty=84; 15'd17458: duty=92; 15'd17459: duty=104; 15'd17460: duty=99; 15'd17461: duty=96; 15'd17462: duty=90; 15'd17463: duty=74;
15'd17464: duty=85; 15'd17465: duty=107; 15'd17466: duty=107; 15'd17467: duty=95; 15'd17468: duty=93; 15'd17469: duty=79; 15'd17470: duty=80; 15'd17471: duty=93;
15'd17472: duty=107; 15'd17473: duty=103; 15'd17474: duty=91; 15'd17475: duty=95; 15'd17476: duty=105; 15'd17477: duty=98; 15'd17478: duty=111; 15'd17479: duty=108;
15'd17480: duty=104; 15'd17481: duty=107; 15'd17482: duty=116; 15'd17483: duty=128; 15'd17484: duty=137; 15'd17485: duty=133; 15'd17486: duty=137; 15'd17487: duty=138;
15'd17488: duty=134; 15'd17489: duty=144; 15'd17490: duty=138; 15'd17491: duty=148; 15'd17492: duty=154; 15'd17493: duty=144; 15'd17494: duty=148; 15'd17495: duty=151;
15'd17496: duty=154; 15'd17497: duty=164; 15'd17498: duty=151; 15'd17499: duty=155; 15'd17500: duty=157; 15'd17501: duty=155; 15'd17502: duty=161; 15'd17503: duty=175;
15'd17504: duty=169; 15'd17505: duty=166; 15'd17506: duty=174; 15'd17507: duty=175; 15'd17508: duty=172; 15'd17509: duty=187; 15'd17510: duty=192; 15'd17511: duty=183;
15'd17512: duty=183; 15'd17513: duty=179; 15'd17514: duty=172; 15'd17515: duty=164; 15'd17516: duty=161; 15'd17517: duty=156; 15'd17518: duty=151; 15'd17519: duty=144;
15'd17520: duty=146; 15'd17521: duty=142; 15'd17522: duty=154; 15'd17523: duty=150; 15'd17524: duty=148; 15'd17525: duty=145; 15'd17526: duty=139; 15'd17527: duty=134;
15'd17528: duty=125; 15'd17529: duty=121; 15'd17530: duty=111; 15'd17531: duty=119; 15'd17532: duty=121; 15'd17533: duty=109; 15'd17534: duty=110; 15'd17535: duty=94;
15'd17536: duty=93; 15'd17537: duty=98; 15'd17538: duty=87; 15'd17539: duty=79; 15'd17540: duty=75; 15'd17541: duty=101; 15'd17542: duty=96; 15'd17543: duty=93;
15'd17544: duty=90; 15'd17545: duty=81; 15'd17546: duty=93; 15'd17547: duty=91; 15'd17548: duty=82; 15'd17549: duty=98; 15'd17550: duty=89; 15'd17551: duty=95;
15'd17552: duty=101; 15'd17553: duty=96; 15'd17554: duty=107; 15'd17555: duty=101; 15'd17556: duty=99; 15'd17557: duty=108; 15'd17558: duty=110; 15'd17559: duty=124;
15'd17560: duty=119; 15'd17561: duty=113; 15'd17562: duty=126; 15'd17563: duty=115; 15'd17564: duty=115; 15'd17565: duty=109; 15'd17566: duty=115; 15'd17567: duty=134;
15'd17568: duty=134; 15'd17569: duty=131; 15'd17570: duty=140; 15'd17571: duty=136; 15'd17572: duty=146; 15'd17573: duty=150; 15'd17574: duty=148; 15'd17575: duty=147;
15'd17576: duty=151; 15'd17577: duty=144; 15'd17578: duty=139; 15'd17579: duty=139; 15'd17580: duty=148; 15'd17581: duty=143; 15'd17582: duty=149; 15'd17583: duty=161;
15'd17584: duty=166; 15'd17585: duty=165; 15'd17586: duty=159; 15'd17587: duty=173; 15'd17588: duty=179; 15'd17589: duty=196; 15'd17590: duty=188; 15'd17591: duty=182;
15'd17592: duty=189; 15'd17593: duty=194; 15'd17594: duty=183; 15'd17595: duty=178; 15'd17596: duty=167; 15'd17597: duty=164; 15'd17598: duty=165; 15'd17599: duty=162;
15'd17600: duty=156; 15'd17601: duty=150; 15'd17602: duty=151; 15'd17603: duty=151; 15'd17604: duty=145; 15'd17605: duty=149; 15'd17606: duty=145; 15'd17607: duty=145;
15'd17608: duty=145; 15'd17609: duty=125; 15'd17610: duty=130; 15'd17611: duty=142; 15'd17612: duty=131; 15'd17613: duty=104; 15'd17614: duty=104; 15'd17615: duty=95;
15'd17616: duty=108; 15'd17617: duty=107; 15'd17618: duty=110; 15'd17619: duty=107; 15'd17620: duty=99; 15'd17621: duty=95; 15'd17622: duty=79; 15'd17623: duty=90;
15'd17624: duty=106; 15'd17625: duty=98; 15'd17626: duty=86; 15'd17627: duty=73; 15'd17628: duty=68; 15'd17629: duty=86; 15'd17630: duty=87; 15'd17631: duty=91;
15'd17632: duty=89; 15'd17633: duty=91; 15'd17634: duty=91; 15'd17635: duty=68; 15'd17636: duty=78; 15'd17637: duty=100; 15'd17638: duty=101; 15'd17639: duty=98;
15'd17640: duty=91; 15'd17641: duty=100; 15'd17642: duty=108; 15'd17643: duty=122; 15'd17644: duty=114; 15'd17645: duty=117; 15'd17646: duty=124; 15'd17647: duty=122;
15'd17648: duty=123; 15'd17649: duty=138; 15'd17650: duty=135; 15'd17651: duty=132; 15'd17652: duty=152; 15'd17653: duty=145; 15'd17654: duty=146; 15'd17655: duty=144;
15'd17656: duty=156; 15'd17657: duty=152; 15'd17658: duty=152; 15'd17659: duty=158; 15'd17660: duty=160; 15'd17661: duty=155; 15'd17662: duty=158; 15'd17663: duty=154;
15'd17664: duty=152; 15'd17665: duty=163; 15'd17666: duty=162; 15'd17667: duty=158; 15'd17668: duty=160; 15'd17669: duty=175; 15'd17670: duty=178; 15'd17671: duty=173;
15'd17672: duty=177; 15'd17673: duty=165; 15'd17674: duty=166; 15'd17675: duty=185; 15'd17676: duty=182; 15'd17677: duty=178; 15'd17678: duty=179; 15'd17679: duty=176;
15'd17680: duty=171; 15'd17681: duty=176; 15'd17682: duty=162; 15'd17683: duty=157; 15'd17684: duty=163; 15'd17685: duty=144; 15'd17686: duty=134; 15'd17687: duty=128;
15'd17688: duty=131; 15'd17689: duty=134; 15'd17690: duty=125; 15'd17691: duty=128; 15'd17692: duty=135; 15'd17693: duty=133; 15'd17694: duty=127; 15'd17695: duty=126;
15'd17696: duty=124; 15'd17697: duty=118; 15'd17698: duty=105; 15'd17699: duty=104; 15'd17700: duty=97; 15'd17701: duty=98; 15'd17702: duty=101; 15'd17703: duty=100;
15'd17704: duty=99; 15'd17705: duty=78; 15'd17706: duty=88; 15'd17707: duty=94; 15'd17708: duty=80; 15'd17709: duty=91; 15'd17710: duty=97; 15'd17711: duty=98;
15'd17712: duty=85; 15'd17713: duty=97; 15'd17714: duty=105; 15'd17715: duty=84; 15'd17716: duty=99; 15'd17717: duty=103; 15'd17718: duty=83; 15'd17719: duty=81;
15'd17720: duty=86; 15'd17721: duty=89; 15'd17722: duty=107; 15'd17723: duty=121; 15'd17724: duty=125; 15'd17725: duty=123; 15'd17726: duty=117; 15'd17727: duty=109;
15'd17728: duty=120; 15'd17729: duty=132; 15'd17730: duty=120; 15'd17731: duty=121; 15'd17732: duty=129; 15'd17733: duty=125; 15'd17734: duty=131; 15'd17735: duty=138;
15'd17736: duty=120; 15'd17737: duty=120; 15'd17738: duty=144; 15'd17739: duty=130; 15'd17740: duty=140; 15'd17741: duty=156; 15'd17742: duty=148; 15'd17743: duty=146;
15'd17744: duty=134; 15'd17745: duty=133; 15'd17746: duty=143; 15'd17747: duty=167; 15'd17748: duty=178; 15'd17749: duty=170; 15'd17750: duty=180; 15'd17751: duty=170;
15'd17752: duty=164; 15'd17753: duty=170; 15'd17754: duty=180; 15'd17755: duty=191; 15'd17756: duty=184; 15'd17757: duty=178; 15'd17758: duty=172; 15'd17759: duty=181;
15'd17760: duty=174; 15'd17761: duty=163; 15'd17762: duty=165; 15'd17763: duty=158; 15'd17764: duty=145; 15'd17765: duty=147; 15'd17766: duty=146; 15'd17767: duty=148;
15'd17768: duty=151; 15'd17769: duty=153; 15'd17770: duty=148; 15'd17771: duty=149; 15'd17772: duty=163; 15'd17773: duty=152; 15'd17774: duty=144; 15'd17775: duty=135;
15'd17776: duty=135; 15'd17777: duty=135; 15'd17778: duty=114; 15'd17779: duty=115; 15'd17780: duty=114; 15'd17781: duty=106; 15'd17782: duty=103; 15'd17783: duty=103;
15'd17784: duty=109; 15'd17785: duty=115; 15'd17786: duty=95; 15'd17787: duty=89; 15'd17788: duty=92; 15'd17789: duty=98; 15'd17790: duty=114; 15'd17791: duty=92;
15'd17792: duty=89; 15'd17793: duty=92; 15'd17794: duty=92; 15'd17795: duty=88; 15'd17796: duty=89; 15'd17797: duty=97; 15'd17798: duty=103; 15'd17799: duty=103;
15'd17800: duty=109; 15'd17801: duty=103; 15'd17802: duty=108; 15'd17803: duty=95; 15'd17804: duty=88; 15'd17805: duty=86; 15'd17806: duty=89; 15'd17807: duty=97;
15'd17808: duty=95; 15'd17809: duty=112; 15'd17810: duty=102; 15'd17811: duty=103; 15'd17812: duty=115; 15'd17813: duty=105; 15'd17814: duty=112; 15'd17815: duty=141;
15'd17816: duty=141; 15'd17817: duty=147; 15'd17818: duty=140; 15'd17819: duty=135; 15'd17820: duty=131; 15'd17821: duty=128; 15'd17822: duty=132; 15'd17823: duty=131;
15'd17824: duty=143; 15'd17825: duty=144; 15'd17826: duty=145; 15'd17827: duty=155; 15'd17828: duty=163; 15'd17829: duty=167; 15'd17830: duty=163; 15'd17831: duty=173;
15'd17832: duty=189; 15'd17833: duty=189; 15'd17834: duty=180; 15'd17835: duty=171; 15'd17836: duty=177; 15'd17837: duty=180; 15'd17838: duty=183; 15'd17839: duty=179;
15'd17840: duty=175; 15'd17841: duty=174; 15'd17842: duty=174; 15'd17843: duty=179; 15'd17844: duty=180; 15'd17845: duty=171; 15'd17846: duty=168; 15'd17847: duty=159;
15'd17848: duty=136; 15'd17849: duty=143; 15'd17850: duty=151; 15'd17851: duty=142; 15'd17852: duty=147; 15'd17853: duty=142; 15'd17854: duty=133; 15'd17855: duty=135;
15'd17856: duty=133; 15'd17857: duty=129; 15'd17858: duty=120; 15'd17859: duty=124; 15'd17860: duty=123; 15'd17861: duty=121; 15'd17862: duty=121; 15'd17863: duty=107;
15'd17864: duty=104; 15'd17865: duty=108; 15'd17866: duty=107; 15'd17867: duty=110; 15'd17868: duty=101; 15'd17869: duty=84; 15'd17870: duty=95; 15'd17871: duty=94;
15'd17872: duty=89; 15'd17873: duty=106; 15'd17874: duty=106; 15'd17875: duty=96; 15'd17876: duty=89; 15'd17877: duty=87; 15'd17878: duty=89; 15'd17879: duty=102;
15'd17880: duty=92; 15'd17881: duty=91; 15'd17882: duty=99; 15'd17883: duty=99; 15'd17884: duty=112; 15'd17885: duty=107; 15'd17886: duty=112; 15'd17887: duty=110;
15'd17888: duty=112; 15'd17889: duty=113; 15'd17890: duty=112; 15'd17891: duty=122; 15'd17892: duty=112; 15'd17893: duty=105; 15'd17894: duty=110; 15'd17895: duty=113;
15'd17896: duty=112; 15'd17897: duty=106; 15'd17898: duty=121; 15'd17899: duty=119; 15'd17900: duty=115; 15'd17901: duty=129; 15'd17902: duty=130; 15'd17903: duty=142;
15'd17904: duty=138; 15'd17905: duty=128; 15'd17906: duty=145; 15'd17907: duty=145; 15'd17908: duty=142; 15'd17909: duty=152; 15'd17910: duty=162; 15'd17911: duty=157;
15'd17912: duty=149; 15'd17913: duty=154; 15'd17914: duty=156; 15'd17915: duty=171; 15'd17916: duty=175; 15'd17917: duty=169; 15'd17918: duty=175; 15'd17919: duty=167;
15'd17920: duty=181; 15'd17921: duty=195; 15'd17922: duty=170; 15'd17923: duty=164; 15'd17924: duty=168; 15'd17925: duty=174; 15'd17926: duty=166; 15'd17927: duty=166;
15'd17928: duty=164; 15'd17929: duty=155; 15'd17930: duty=153; 15'd17931: duty=152; 15'd17932: duty=155; 15'd17933: duty=155; 15'd17934: duty=161; 15'd17935: duty=155;
15'd17936: duty=149; 15'd17937: duty=151; 15'd17938: duty=139; 15'd17939: duty=138; 15'd17940: duty=128; 15'd17941: duty=124; 15'd17942: duty=133; 15'd17943: duty=129;
15'd17944: duty=134; 15'd17945: duty=119; 15'd17946: duty=116; 15'd17947: duty=119; 15'd17948: duty=119; 15'd17949: duty=118; 15'd17950: duty=114; 15'd17951: duty=107;
15'd17952: duty=104; 15'd17953: duty=101; 15'd17954: duty=94; 15'd17955: duty=95; 15'd17956: duty=93; 15'd17957: duty=95; 15'd17958: duty=90; 15'd17959: duty=86;
15'd17960: duty=96; 15'd17961: duty=101; 15'd17962: duty=101; 15'd17963: duty=101; 15'd17964: duty=104; 15'd17965: duty=98; 15'd17966: duty=108; 15'd17967: duty=112;
15'd17968: duty=88; 15'd17969: duty=81; 15'd17970: duty=90; 15'd17971: duty=108; 15'd17972: duty=109; 15'd17973: duty=92; 15'd17974: duty=91; 15'd17975: duty=96;
15'd17976: duty=103; 15'd17977: duty=111; 15'd17978: duty=115; 15'd17979: duty=126; 15'd17980: duty=121; 15'd17981: duty=127; 15'd17982: duty=132; 15'd17983: duty=121;
15'd17984: duty=134; 15'd17985: duty=133; 15'd17986: duty=116; 15'd17987: duty=122; 15'd17988: duty=127; 15'd17989: duty=133; 15'd17990: duty=143; 15'd17991: duty=136;
15'd17992: duty=132; 15'd17993: duty=140; 15'd17994: duty=140; 15'd17995: duty=149; 15'd17996: duty=165; 15'd17997: duty=170; 15'd17998: duty=159; 15'd17999: duty=171;
15'd18000: duty=176; 15'd18001: duty=171; 15'd18002: duty=194; 15'd18003: duty=195; 15'd18004: duty=183; 15'd18005: duty=182; 15'd18006: duty=183; 15'd18007: duty=183;
15'd18008: duty=179; 15'd18009: duty=168; 15'd18010: duty=171; 15'd18011: duty=174; 15'd18012: duty=160; 15'd18013: duty=159; 15'd18014: duty=157; 15'd18015: duty=158;
15'd18016: duty=152; 15'd18017: duty=145; 15'd18018: duty=151; 15'd18019: duty=152; 15'd18020: duty=155; 15'd18021: duty=147; 15'd18022: duty=137; 15'd18023: duty=147;
15'd18024: duty=141; 15'd18025: duty=126; 15'd18026: duty=127; 15'd18027: duty=112; 15'd18028: duty=113; 15'd18029: duty=104; 15'd18030: duty=103; 15'd18031: duty=109;
15'd18032: duty=108; 15'd18033: duty=103; 15'd18034: duty=88; 15'd18035: duty=89; 15'd18036: duty=105; 15'd18037: duty=111; 15'd18038: duty=103; 15'd18039: duty=104;
15'd18040: duty=99; 15'd18041: duty=90; 15'd18042: duty=85; 15'd18043: duty=91; 15'd18044: duty=91; 15'd18045: duty=83; 15'd18046: duty=92; 15'd18047: duty=93;
15'd18048: duty=100; 15'd18049: duty=100; 15'd18050: duty=101; 15'd18051: duty=118; 15'd18052: duty=108; 15'd18053: duty=107; 15'd18054: duty=102; 15'd18055: duty=106;
15'd18056: duty=117; 15'd18057: duty=123; 15'd18058: duty=112; 15'd18059: duty=107; 15'd18060: duty=107; 15'd18061: duty=119; 15'd18062: duty=124; 15'd18063: duty=113;
15'd18064: duty=115; 15'd18065: duty=127; 15'd18066: duty=140; 15'd18067: duty=134; 15'd18068: duty=138; 15'd18069: duty=145; 15'd18070: duty=136; 15'd18071: duty=131;
15'd18072: duty=142; 15'd18073: duty=137; 15'd18074: duty=142; 15'd18075: duty=140; 15'd18076: duty=150; 15'd18077: duty=157; 15'd18078: duty=158; 15'd18079: duty=157;
15'd18080: duty=156; 15'd18081: duty=159; 15'd18082: duty=167; 15'd18083: duty=175; 15'd18084: duty=173; 15'd18085: duty=168; 15'd18086: duty=168; 15'd18087: duty=179;
15'd18088: duty=168; 15'd18089: duty=169; 15'd18090: duty=171; 15'd18091: duty=166; 15'd18092: duty=161; 15'd18093: duty=154; 15'd18094: duty=154; 15'd18095: duty=152;
15'd18096: duty=148; 15'd18097: duty=151; 15'd18098: duty=145; 15'd18099: duty=148; 15'd18100: duty=153; 15'd18101: duty=148; 15'd18102: duty=147; 15'd18103: duty=134;
15'd18104: duty=131; 15'd18105: duty=141; 15'd18106: duty=131; 15'd18107: duty=128; 15'd18108: duty=123; 15'd18109: duty=119; 15'd18110: duty=122; 15'd18111: duty=125;
15'd18112: duty=127; 15'd18113: duty=113; 15'd18114: duty=106; 15'd18115: duty=104; 15'd18116: duty=102; 15'd18117: duty=104; 15'd18118: duty=104; 15'd18119: duty=102;
15'd18120: duty=102; 15'd18121: duty=98; 15'd18122: duty=99; 15'd18123: duty=109; 15'd18124: duty=102; 15'd18125: duty=95; 15'd18126: duty=99; 15'd18127: duty=87;
15'd18128: duty=88; 15'd18129: duty=101; 15'd18130: duty=96; 15'd18131: duty=87; 15'd18132: duty=102; 15'd18133: duty=101; 15'd18134: duty=105; 15'd18135: duty=115;
15'd18136: duty=125; 15'd18137: duty=121; 15'd18138: duty=120; 15'd18139: duty=115; 15'd18140: duty=104; 15'd18141: duty=113; 15'd18142: duty=122; 15'd18143: duty=127;
15'd18144: duty=125; 15'd18145: duty=132; 15'd18146: duty=128; 15'd18147: duty=133; 15'd18148: duty=132; 15'd18149: duty=136; 15'd18150: duty=158; 15'd18151: duty=159;
15'd18152: duty=141; 15'd18153: duty=149; 15'd18154: duty=141; 15'd18155: duty=153; 15'd18156: duty=159; 15'd18157: duty=149; 15'd18158: duty=151; 15'd18159: duty=162;
15'd18160: duty=169; 15'd18161: duty=161; 15'd18162: duty=160; 15'd18163: duty=166; 15'd18164: duty=163; 15'd18165: duty=165; 15'd18166: duty=175; 15'd18167: duty=177;
15'd18168: duty=178; 15'd18169: duty=166; 15'd18170: duty=173; 15'd18171: duty=173; 15'd18172: duty=169; 15'd18173: duty=165; 15'd18174: duty=162; 15'd18175: duty=147;
15'd18176: duty=147; 15'd18177: duty=139; 15'd18178: duty=143; 15'd18179: duty=144; 15'd18180: duty=137; 15'd18181: duty=134; 15'd18182: duty=132; 15'd18183: duty=126;
15'd18184: duty=117; 15'd18185: duty=126; 15'd18186: duty=136; 15'd18187: duty=123; 15'd18188: duty=129; 15'd18189: duty=124; 15'd18190: duty=120; 15'd18191: duty=124;
15'd18192: duty=114; 15'd18193: duty=115; 15'd18194: duty=114; 15'd18195: duty=107; 15'd18196: duty=102; 15'd18197: duty=104; 15'd18198: duty=94; 15'd18199: duty=92;
15'd18200: duty=86; 15'd18201: duty=93; 15'd18202: duty=94; 15'd18203: duty=100; 15'd18204: duty=108; 15'd18205: duty=98; 15'd18206: duty=85; 15'd18207: duty=78;
15'd18208: duty=81; 15'd18209: duty=97; 15'd18210: duty=102; 15'd18211: duty=107; 15'd18212: duty=103; 15'd18213: duty=109; 15'd18214: duty=118; 15'd18215: duty=120;
15'd18216: duty=116; 15'd18217: duty=112; 15'd18218: duty=108; 15'd18219: duty=109; 15'd18220: duty=106; 15'd18221: duty=101; 15'd18222: duty=125; 15'd18223: duty=113;
15'd18224: duty=105; 15'd18225: duty=105; 15'd18226: duty=116; 15'd18227: duty=131; 15'd18228: duty=135; 15'd18229: duty=142; 15'd18230: duty=149; 15'd18231: duty=148;
15'd18232: duty=139; 15'd18233: duty=147; 15'd18234: duty=143; 15'd18235: duty=140; 15'd18236: duty=145; 15'd18237: duty=154; 15'd18238: duty=162; 15'd18239: duty=177;
15'd18240: duty=164; 15'd18241: duty=160; 15'd18242: duty=180; 15'd18243: duty=166; 15'd18244: duty=170; 15'd18245: duty=181; 15'd18246: duty=185; 15'd18247: duty=185;
15'd18248: duty=178; 15'd18249: duty=179; 15'd18250: duty=180; 15'd18251: duty=179; 15'd18252: duty=185; 15'd18253: duty=169; 15'd18254: duty=161; 15'd18255: duty=157;
15'd18256: duty=150; 15'd18257: duty=145; 15'd18258: duty=147; 15'd18259: duty=141; 15'd18260: duty=142; 15'd18261: duty=145; 15'd18262: duty=139; 15'd18263: duty=141;
15'd18264: duty=142; 15'd18265: duty=131; 15'd18266: duty=134; 15'd18267: duty=131; 15'd18268: duty=123; 15'd18269: duty=129; 15'd18270: duty=115; 15'd18271: duty=104;
15'd18272: duty=105; 15'd18273: duty=110; 15'd18274: duty=100; 15'd18275: duty=101; 15'd18276: duty=109; 15'd18277: duty=100; 15'd18278: duty=98; 15'd18279: duty=102;
15'd18280: duty=81; 15'd18281: duty=91; 15'd18282: duty=91; 15'd18283: duty=73; 15'd18284: duty=77; 15'd18285: duty=105; 15'd18286: duty=108; 15'd18287: duty=96;
15'd18288: duty=94; 15'd18289: duty=93; 15'd18290: duty=89; 15'd18291: duty=97; 15'd18292: duty=106; 15'd18293: duty=117; 15'd18294: duty=117; 15'd18295: duty=91;
15'd18296: duty=101; 15'd18297: duty=117; 15'd18298: duty=120; 15'd18299: duty=120; 15'd18300: duty=123; 15'd18301: duty=119; 15'd18302: duty=125; 15'd18303: duty=132;
15'd18304: duty=146; 15'd18305: duty=136; 15'd18306: duty=142; 15'd18307: duty=142; 15'd18308: duty=136; 15'd18309: duty=147; 15'd18310: duty=150; 15'd18311: duty=147;
15'd18312: duty=141; 15'd18313: duty=128; 15'd18314: duty=132; 15'd18315: duty=150; 15'd18316: duty=159; 15'd18317: duty=152; 15'd18318: duty=150; 15'd18319: duty=155;
15'd18320: duty=156; 15'd18321: duty=161; 15'd18322: duty=159; 15'd18323: duty=152; 15'd18324: duty=166; 15'd18325: duty=174; 15'd18326: duty=161; 15'd18327: duty=162;
15'd18328: duty=164; 15'd18329: duty=174; 15'd18330: duty=170; 15'd18331: duty=168; 15'd18332: duty=168; 15'd18333: duty=171; 15'd18334: duty=173; 15'd18335: duty=160;
15'd18336: duty=150; 15'd18337: duty=145; 15'd18338: duty=137; 15'd18339: duty=148; 15'd18340: duty=132; 15'd18341: duty=128; 15'd18342: duty=138; 15'd18343: duty=134;
15'd18344: duty=128; 15'd18345: duty=127; 15'd18346: duty=122; 15'd18347: duty=124; 15'd18348: duty=134; 15'd18349: duty=133; 15'd18350: duty=127; 15'd18351: duty=122;
15'd18352: duty=135; 15'd18353: duty=117; 15'd18354: duty=110; 15'd18355: duty=112; 15'd18356: duty=105; 15'd18357: duty=101; 15'd18358: duty=101; 15'd18359: duty=92;
15'd18360: duty=94; 15'd18361: duty=100; 15'd18362: duty=104; 15'd18363: duty=92; 15'd18364: duty=99; 15'd18365: duty=110; 15'd18366: duty=90; 15'd18367: duty=89;
15'd18368: duty=101; 15'd18369: duty=101; 15'd18370: duty=104; 15'd18371: duty=96; 15'd18372: duty=107; 15'd18373: duty=107; 15'd18374: duty=93; 15'd18375: duty=105;
15'd18376: duty=105; 15'd18377: duty=113; 15'd18378: duty=124; 15'd18379: duty=118; 15'd18380: duty=113; 15'd18381: duty=118; 15'd18382: duty=119; 15'd18383: duty=127;
15'd18384: duty=126; 15'd18385: duty=121; 15'd18386: duty=118; 15'd18387: duty=128; 15'd18388: duty=131; 15'd18389: duty=119; 15'd18390: duty=124; 15'd18391: duty=145;
15'd18392: duty=138; 15'd18393: duty=131; 15'd18394: duty=134; 15'd18395: duty=142; 15'd18396: duty=159; 15'd18397: duty=140; 15'd18398: duty=139; 15'd18399: duty=148;
15'd18400: duty=160; 15'd18401: duty=160; 15'd18402: duty=167; 15'd18403: duty=163; 15'd18404: duty=150; 15'd18405: duty=157; 15'd18406: duty=159; 15'd18407: duty=171;
15'd18408: duty=175; 15'd18409: duty=176; 15'd18410: duty=170; 15'd18411: duty=171; 15'd18412: duty=176; 15'd18413: duty=177; 15'd18414: duty=169; 15'd18415: duty=157;
15'd18416: duty=156; 15'd18417: duty=162; 15'd18418: duty=164; 15'd18419: duty=153; 15'd18420: duty=154; 15'd18421: duty=152; 15'd18422: duty=150; 15'd18423: duty=148;
15'd18424: duty=142; 15'd18425: duty=142; 15'd18426: duty=142; 15'd18427: duty=134; 15'd18428: duty=129; 15'd18429: duty=124; 15'd18430: duty=131; 15'd18431: duty=127;
15'd18432: duty=117; 15'd18433: duty=122; 15'd18434: duty=117; 15'd18435: duty=119; 15'd18436: duty=118; 15'd18437: duty=128; 15'd18438: duty=124; 15'd18439: duty=105;
15'd18440: duty=100; 15'd18441: duty=105; 15'd18442: duty=106; 15'd18443: duty=111; 15'd18444: duty=97; 15'd18445: duty=91; 15'd18446: duty=105; 15'd18447: duty=105;
15'd18448: duty=104; 15'd18449: duty=96; 15'd18450: duty=89; 15'd18451: duty=85; 15'd18452: duty=89; 15'd18453: duty=88; 15'd18454: duty=100; 15'd18455: duty=103;
15'd18456: duty=106; 15'd18457: duty=97; 15'd18458: duty=98; 15'd18459: duty=110; 15'd18460: duty=115; 15'd18461: duty=117; 15'd18462: duty=101; 15'd18463: duty=100;
15'd18464: duty=114; 15'd18465: duty=119; 15'd18466: duty=124; 15'd18467: duty=127; 15'd18468: duty=118; 15'd18469: duty=124; 15'd18470: duty=127; 15'd18471: duty=132;
15'd18472: duty=136; 15'd18473: duty=134; 15'd18474: duty=136; 15'd18475: duty=133; 15'd18476: duty=143; 15'd18477: duty=148; 15'd18478: duty=151; 15'd18479: duty=154;
15'd18480: duty=142; 15'd18481: duty=151; 15'd18482: duty=153; 15'd18483: duty=158; 15'd18484: duty=165; 15'd18485: duty=158; 15'd18486: duty=150; 15'd18487: duty=151;
15'd18488: duty=161; 15'd18489: duty=169; 15'd18490: duty=176; 15'd18491: duty=175; 15'd18492: duty=175; 15'd18493: duty=174; 15'd18494: duty=180; 15'd18495: duty=179;
15'd18496: duty=179; 15'd18497: duty=169; 15'd18498: duty=158; 15'd18499: duty=161; 15'd18500: duty=158; 15'd18501: duty=152; 15'd18502: duty=146; 15'd18503: duty=140;
15'd18504: duty=139; 15'd18505: duty=140; 15'd18506: duty=149; 15'd18507: duty=144; 15'd18508: duty=147; 15'd18509: duty=142; 15'd18510: duty=127; 15'd18511: duty=130;
15'd18512: duty=121; 15'd18513: duty=119; 15'd18514: duty=126; 15'd18515: duty=111; 15'd18516: duty=104; 15'd18517: duty=115; 15'd18518: duty=107; 15'd18519: duty=99;
15'd18520: duty=103; 15'd18521: duty=111; 15'd18522: duty=112; 15'd18523: duty=99; 15'd18524: duty=87; 15'd18525: duty=99; 15'd18526: duty=94; 15'd18527: duty=88;
15'd18528: duty=93; 15'd18529: duty=101; 15'd18530: duty=94; 15'd18531: duty=96; 15'd18532: duty=102; 15'd18533: duty=102; 15'd18534: duty=107; 15'd18535: duty=102;
15'd18536: duty=103; 15'd18537: duty=106; 15'd18538: duty=107; 15'd18539: duty=107; 15'd18540: duty=108; 15'd18541: duty=101; 15'd18542: duty=119; 15'd18543: duty=117;
15'd18544: duty=119; 15'd18545: duty=130; 15'd18546: duty=122; 15'd18547: duty=98; 15'd18548: duty=105; 15'd18549: duty=126; 15'd18550: duty=131; 15'd18551: duty=136;
15'd18552: duty=135; 15'd18553: duty=141; 15'd18554: duty=134; 15'd18555: duty=133; 15'd18556: duty=142; 15'd18557: duty=134; 15'd18558: duty=140; 15'd18559: duty=133;
15'd18560: duty=136; 15'd18561: duty=160; 15'd18562: duty=143; 15'd18563: duty=148; 15'd18564: duty=144; 15'd18565: duty=137; 15'd18566: duty=160; 15'd18567: duty=177;
15'd18568: duty=173; 15'd18569: duty=181; 15'd18570: duty=188; 15'd18571: duty=185; 15'd18572: duty=181; 15'd18573: duty=180; 15'd18574: duty=182; 15'd18575: duty=174;
15'd18576: duty=169; 15'd18577: duty=163; 15'd18578: duty=170; 15'd18579: duty=165; 15'd18580: duty=161; 15'd18581: duty=157; 15'd18582: duty=153; 15'd18583: duty=160;
15'd18584: duty=167; 15'd18585: duty=169; 15'd18586: duty=165; 15'd18587: duty=150; 15'd18588: duty=153; 15'd18589: duty=155; 15'd18590: duty=143; 15'd18591: duty=139;
15'd18592: duty=126; 15'd18593: duty=108; 15'd18594: duty=106; 15'd18595: duty=113; 15'd18596: duty=115; 15'd18597: duty=106; 15'd18598: duty=108; 15'd18599: duty=94;
15'd18600: duty=91; 15'd18601: duty=108; 15'd18602: duty=93; 15'd18603: duty=103; 15'd18604: duty=94; 15'd18605: duty=82; 15'd18606: duty=94; 15'd18607: duty=105;
15'd18608: duty=78; 15'd18609: duty=63; 15'd18610: duty=80; 15'd18611: duty=88; 15'd18612: duty=90; 15'd18613: duty=82; 15'd18614: duty=104; 15'd18615: duty=111;
15'd18616: duty=109; 15'd18617: duty=105; 15'd18618: duty=114; 15'd18619: duty=117; 15'd18620: duty=92; 15'd18621: duty=91; 15'd18622: duty=99; 15'd18623: duty=97;
15'd18624: duty=112; 15'd18625: duty=108; 15'd18626: duty=95; 15'd18627: duty=117; 15'd18628: duty=118; 15'd18629: duty=122; 15'd18630: duty=126; 15'd18631: duty=128;
15'd18632: duty=130; 15'd18633: duty=134; 15'd18634: duty=155; 15'd18635: duty=142; 15'd18636: duty=146; 15'd18637: duty=154; 15'd18638: duty=139; 15'd18639: duty=146;
15'd18640: duty=156; 15'd18641: duty=160; 15'd18642: duty=159; 15'd18643: duty=151; 15'd18644: duty=153; 15'd18645: duty=157; 15'd18646: duty=161; 15'd18647: duty=170;
15'd18648: duty=159; 15'd18649: duty=170; 15'd18650: duty=180; 15'd18651: duty=168; 15'd18652: duty=176; 15'd18653: duty=194; 15'd18654: duty=189; 15'd18655: duty=179;
15'd18656: duty=180; 15'd18657: duty=174; 15'd18658: duty=179; 15'd18659: duty=182; 15'd18660: duty=168; 15'd18661: duty=162; 15'd18662: duty=156; 15'd18663: duty=150;
15'd18664: duty=144; 15'd18665: duty=146; 15'd18666: duty=151; 15'd18667: duty=146; 15'd18668: duty=135; 15'd18669: duty=128; 15'd18670: duty=132; 15'd18671: duty=128;
15'd18672: duty=127; 15'd18673: duty=121; 15'd18674: duty=120; 15'd18675: duty=120; 15'd18676: duty=119; 15'd18677: duty=118; 15'd18678: duty=107; 15'd18679: duty=110;
15'd18680: duty=108; 15'd18681: duty=96; 15'd18682: duty=97; 15'd18683: duty=115; 15'd18684: duty=94; 15'd18685: duty=82; 15'd18686: duty=98; 15'd18687: duty=89;
15'd18688: duty=86; 15'd18689: duty=83; 15'd18690: duty=97; 15'd18691: duty=96; 15'd18692: duty=85; 15'd18693: duty=86; 15'd18694: duty=87; 15'd18695: duty=78;
15'd18696: duty=90; 15'd18697: duty=104; 15'd18698: duty=88; 15'd18699: duty=98; 15'd18700: duty=97; 15'd18701: duty=100; 15'd18702: duty=108; 15'd18703: duty=112;
15'd18704: duty=115; 15'd18705: duty=115; 15'd18706: duty=124; 15'd18707: duty=112; 15'd18708: duty=120; 15'd18709: duty=125; 15'd18710: duty=119; 15'd18711: duty=133;
15'd18712: duty=145; 15'd18713: duty=139; 15'd18714: duty=132; 15'd18715: duty=141; 15'd18716: duty=149; 15'd18717: duty=149; 15'd18718: duty=155; 15'd18719: duty=156;
15'd18720: duty=143; 15'd18721: duty=144; 15'd18722: duty=145; 15'd18723: duty=153; 15'd18724: duty=165; 15'd18725: duty=160; 15'd18726: duty=157; 15'd18727: duty=152;
15'd18728: duty=154; 15'd18729: duty=167; 15'd18730: duty=170; 15'd18731: duty=178; 15'd18732: duty=175; 15'd18733: duty=172; 15'd18734: duty=177; 15'd18735: duty=182;
15'd18736: duty=178; 15'd18737: duty=179; 15'd18738: duty=177; 15'd18739: duty=173; 15'd18740: duty=170; 15'd18741: duty=168; 15'd18742: duty=169; 15'd18743: duty=154;
15'd18744: duty=149; 15'd18745: duty=151; 15'd18746: duty=152; 15'd18747: duty=151; 15'd18748: duty=154; 15'd18749: duty=145; 15'd18750: duty=146; 15'd18751: duty=149;
15'd18752: duty=137; 15'd18753: duty=138; 15'd18754: duty=127; 15'd18755: duty=115; 15'd18756: duty=121; 15'd18757: duty=126; 15'd18758: duty=128; 15'd18759: duty=113;
15'd18760: duty=117; 15'd18761: duty=112; 15'd18762: duty=90; 15'd18763: duty=93; 15'd18764: duty=104; 15'd18765: duty=95; 15'd18766: duty=98; 15'd18767: duty=93;
15'd18768: duty=76; 15'd18769: duty=84; 15'd18770: duty=84; 15'd18771: duty=82; 15'd18772: duty=82; 15'd18773: duty=86; 15'd18774: duty=74; 15'd18775: duty=69;
15'd18776: duty=85; 15'd18777: duty=98; 15'd18778: duty=84; 15'd18779: duty=83; 15'd18780: duty=87; 15'd18781: duty=92; 15'd18782: duty=108; 15'd18783: duty=103;
15'd18784: duty=110; 15'd18785: duty=116; 15'd18786: duty=110; 15'd18787: duty=110; 15'd18788: duty=121; 15'd18789: duty=116; 15'd18790: duty=117; 15'd18791: duty=110;
15'd18792: duty=104; 15'd18793: duty=120; 15'd18794: duty=113; 15'd18795: duty=129; 15'd18796: duty=145; 15'd18797: duty=135; 15'd18798: duty=141; 15'd18799: duty=142;
15'd18800: duty=141; 15'd18801: duty=165; 15'd18802: duty=161; 15'd18803: duty=156; 15'd18804: duty=154; 15'd18805: duty=150; 15'd18806: duty=154; 15'd18807: duty=162;
15'd18808: duty=171; 15'd18809: duty=161; 15'd18810: duty=171; 15'd18811: duty=182; 15'd18812: duty=183; 15'd18813: duty=182; 15'd18814: duty=183; 15'd18815: duty=181;
15'd18816: duty=183; 15'd18817: duty=196; 15'd18818: duty=188; 15'd18819: duty=184; 15'd18820: duty=181; 15'd18821: duty=167; 15'd18822: duty=177; 15'd18823: duty=176;
15'd18824: duty=166; 15'd18825: duty=156; 15'd18826: duty=160; 15'd18827: duty=165; 15'd18828: duty=158; 15'd18829: duty=155; 15'd18830: duty=154; 15'd18831: duty=154;
15'd18832: duty=148; 15'd18833: duty=142; 15'd18834: duty=134; 15'd18835: duty=131; 15'd18836: duty=129; 15'd18837: duty=118; 15'd18838: duty=121; 15'd18839: duty=110;
15'd18840: duty=102; 15'd18841: duty=107; 15'd18842: duty=117; 15'd18843: duty=118; 15'd18844: duty=98; 15'd18845: duty=106; 15'd18846: duty=99; 15'd18847: duty=86;
15'd18848: duty=79; 15'd18849: duty=86; 15'd18850: duty=99; 15'd18851: duty=92; 15'd18852: duty=88; 15'd18853: duty=95; 15'd18854: duty=105; 15'd18855: duty=107;
15'd18856: duty=94; 15'd18857: duty=79; 15'd18858: duty=84; 15'd18859: duty=93; 15'd18860: duty=90; 15'd18861: duty=98; 15'd18862: duty=93; 15'd18863: duty=87;
15'd18864: duty=94; 15'd18865: duty=97; 15'd18866: duty=93; 15'd18867: duty=93; 15'd18868: duty=104; 15'd18869: duty=103; 15'd18870: duty=117; 15'd18871: duty=120;
15'd18872: duty=110; 15'd18873: duty=108; 15'd18874: duty=102; 15'd18875: duty=101; 15'd18876: duty=116; 15'd18877: duty=120; 15'd18878: duty=119; 15'd18879: duty=126;
15'd18880: duty=129; 15'd18881: duty=133; 15'd18882: duty=149; 15'd18883: duty=154; 15'd18884: duty=143; 15'd18885: duty=145; 15'd18886: duty=151; 15'd18887: duty=152;
15'd18888: duty=166; 15'd18889: duty=170; 15'd18890: duty=176; 15'd18891: duty=171; 15'd18892: duty=170; 15'd18893: duty=167; 15'd18894: duty=169; 15'd18895: duty=191;
15'd18896: duty=188; 15'd18897: duty=179; 15'd18898: duty=175; 15'd18899: duty=184; 15'd18900: duty=180; 15'd18901: duty=177; 15'd18902: duty=165; 15'd18903: duty=156;
15'd18904: duty=160; 15'd18905: duty=164; 15'd18906: duty=173; 15'd18907: duty=178; 15'd18908: duty=164; 15'd18909: duty=159; 15'd18910: duty=157; 15'd18911: duty=151;
15'd18912: duty=156; 15'd18913: duty=162; 15'd18914: duty=159; 15'd18915: duty=146; 15'd18916: duty=134; 15'd18917: duty=134; 15'd18918: duty=145; 15'd18919: duty=142;
15'd18920: duty=135; 15'd18921: duty=127; 15'd18922: duty=121; 15'd18923: duty=127; 15'd18924: duty=127; 15'd18925: duty=109; 15'd18926: duty=98; 15'd18927: duty=100;
15'd18928: duty=112; 15'd18929: duty=110; 15'd18930: duty=99; 15'd18931: duty=97; 15'd18932: duty=99; 15'd18933: duty=91; 15'd18934: duty=81; 15'd18935: duty=85;
15'd18936: duty=87; 15'd18937: duty=84; 15'd18938: duty=78; 15'd18939: duty=76; 15'd18940: duty=83; 15'd18941: duty=73; 15'd18942: duty=64; 15'd18943: duty=73;
15'd18944: duty=82; 15'd18945: duty=94; 15'd18946: duty=100; 15'd18947: duty=96; 15'd18948: duty=86; 15'd18949: duty=90; 15'd18950: duty=105; 15'd18951: duty=113;
15'd18952: duty=102; 15'd18953: duty=117; 15'd18954: duty=107; 15'd18955: duty=106; 15'd18956: duty=128; 15'd18957: duty=129; 15'd18958: duty=131; 15'd18959: duty=121;
15'd18960: duty=128; 15'd18961: duty=138; 15'd18962: duty=146; 15'd18963: duty=142; 15'd18964: duty=138; 15'd18965: duty=139; 15'd18966: duty=145; 15'd18967: duty=151;
15'd18968: duty=154; 15'd18969: duty=156; 15'd18970: duty=155; 15'd18971: duty=162; 15'd18972: duty=162; 15'd18973: duty=167; 15'd18974: duty=179; 15'd18975: duty=188;
15'd18976: duty=191; 15'd18977: duty=193; 15'd18978: duty=189; 15'd18979: duty=186; 15'd18980: duty=187; 15'd18981: duty=173; 15'd18982: duty=171; 15'd18983: duty=168;
15'd18984: duty=168; 15'd18985: duty=172; 15'd18986: duty=171; 15'd18987: duty=163; 15'd18988: duty=154; 15'd18989: duty=157; 15'd18990: duty=159; 15'd18991: duty=149;
15'd18992: duty=148; 15'd18993: duty=157; 15'd18994: duty=149; 15'd18995: duty=142; 15'd18996: duty=134; 15'd18997: duty=132; 15'd18998: duty=129; 15'd18999: duty=119;
15'd19000: duty=119; 15'd19001: duty=118; 15'd19002: duty=118; 15'd19003: duty=123; 15'd19004: duty=116; 15'd19005: duty=105; 15'd19006: duty=101; 15'd19007: duty=105;
15'd19008: duty=105; 15'd19009: duty=107; 15'd19010: duty=99; 15'd19011: duty=104; 15'd19012: duty=113; 15'd19013: duty=92; 15'd19014: duty=78; 15'd19015: duty=92;
15'd19016: duty=107; 15'd19017: duty=105; 15'd19018: duty=94; 15'd19019: duty=96; 15'd19020: duty=96; 15'd19021: duty=97; 15'd19022: duty=99; 15'd19023: duty=82;
15'd19024: duty=81; 15'd19025: duty=84; 15'd19026: duty=93; 15'd19027: duty=90; 15'd19028: duty=99; 15'd19029: duty=101; 15'd19030: duty=108; 15'd19031: duty=110;
15'd19032: duty=108; 15'd19033: duty=117; 15'd19034: duty=124; 15'd19035: duty=124; 15'd19036: duty=110; 15'd19037: duty=128; 15'd19038: duty=136; 15'd19039: duty=145;
15'd19040: duty=134; 15'd19041: duty=129; 15'd19042: duty=126; 15'd19043: duty=133; 15'd19044: duty=137; 15'd19045: duty=128; 15'd19046: duty=137; 15'd19047: duty=145;
15'd19048: duty=159; 15'd19049: duty=150; 15'd19050: duty=154; 15'd19051: duty=159; 15'd19052: duty=168; 15'd19053: duty=170; 15'd19054: duty=173; 15'd19055: duty=186;
15'd19056: duty=199; 15'd19057: duty=197; 15'd19058: duty=185; 15'd19059: duty=183; 15'd19060: duty=185; 15'd19061: duty=176; 15'd19062: duty=164; 15'd19063: duty=162;
15'd19064: duty=171; 15'd19065: duty=180; 15'd19066: duty=171; 15'd19067: duty=168; 15'd19068: duty=162; 15'd19069: duty=162; 15'd19070: duty=155; 15'd19071: duty=149;
15'd19072: duty=158; 15'd19073: duty=160; 15'd19074: duty=144; 15'd19075: duty=137; 15'd19076: duty=131; 15'd19077: duty=129; 15'd19078: duty=124; 15'd19079: duty=121;
15'd19080: duty=131; 15'd19081: duty=129; 15'd19082: duty=119; 15'd19083: duty=104; 15'd19084: duty=119; 15'd19085: duty=119; 15'd19086: duty=110; 15'd19087: duty=115;
15'd19088: duty=106; 15'd19089: duty=94; 15'd19090: duty=102; 15'd19091: duty=91; 15'd19092: duty=95; 15'd19093: duty=104; 15'd19094: duty=89; 15'd19095: duty=95;
15'd19096: duty=88; 15'd19097: duty=95; 15'd19098: duty=98; 15'd19099: duty=88; 15'd19100: duty=101; 15'd19101: duty=95; 15'd19102: duty=85; 15'd19103: duty=96;
15'd19104: duty=85; 15'd19105: duty=81; 15'd19106: duty=90; 15'd19107: duty=91; 15'd19108: duty=93; 15'd19109: duty=99; 15'd19110: duty=102; 15'd19111: duty=113;
15'd19112: duty=114; 15'd19113: duty=108; 15'd19114: duty=118; 15'd19115: duty=112; 15'd19116: duty=110; 15'd19117: duty=124; 15'd19118: duty=115; 15'd19119: duty=104;
15'd19120: duty=116; 15'd19121: duty=131; 15'd19122: duty=134; 15'd19123: duty=144; 15'd19124: duty=140; 15'd19125: duty=147; 15'd19126: duty=150; 15'd19127: duty=151;
15'd19128: duty=157; 15'd19129: duty=141; 15'd19130: duty=163; 15'd19131: duty=162; 15'd19132: duty=168; 15'd19133: duty=174; 15'd19134: duty=162; 15'd19135: duty=173;
15'd19136: duty=186; 15'd19137: duty=187; 15'd19138: duty=179; 15'd19139: duty=196; 15'd19140: duty=202; 15'd19141: duty=190; 15'd19142: duty=183; 15'd19143: duty=173;
15'd19144: duty=160; 15'd19145: duty=160; 15'd19146: duty=173; 15'd19147: duty=171; 15'd19148: duty=168; 15'd19149: duty=157; 15'd19150: duty=148; 15'd19151: duty=150;
15'd19152: duty=152; 15'd19153: duty=144; 15'd19154: duty=148; 15'd19155: duty=153; 15'd19156: duty=146; 15'd19157: duty=140; 15'd19158: duty=124; 15'd19159: duty=124;
15'd19160: duty=122; 15'd19161: duty=119; 15'd19162: duty=117; 15'd19163: duty=109; 15'd19164: duty=107; 15'd19165: duty=116; 15'd19166: duty=119; 15'd19167: duty=116;
15'd19168: duty=117; 15'd19169: duty=113; 15'd19170: duty=96; 15'd19171: duty=96; 15'd19172: duty=105; 15'd19173: duty=101; 15'd19174: duty=99; 15'd19175: duty=92;
15'd19176: duty=88; 15'd19177: duty=101; 15'd19178: duty=99; 15'd19179: duty=112; 15'd19180: duty=92; 15'd19181: duty=81; 15'd19182: duty=96; 15'd19183: duty=92;
15'd19184: duty=96; 15'd19185: duty=93; 15'd19186: duty=99; 15'd19187: duty=93; 15'd19188: duty=95; 15'd19189: duty=105; 15'd19190: duty=118; 15'd19191: duty=113;
15'd19192: duty=118; 15'd19193: duty=118; 15'd19194: duty=107; 15'd19195: duty=118; 15'd19196: duty=109; 15'd19197: duty=107; 15'd19198: duty=106; 15'd19199: duty=107;
15'd19200: duty=113; 15'd19201: duty=113; 15'd19202: duty=121; 15'd19203: duty=135; 15'd19204: duty=142; 15'd19205: duty=143; 15'd19206: duty=130; 15'd19207: duty=129;
15'd19208: duty=144; 15'd19209: duty=140; 15'd19210: duty=144; 15'd19211: duty=155; 15'd19212: duty=149; 15'd19213: duty=154; 15'd19214: duty=161; 15'd19215: duty=161;
15'd19216: duty=178; 15'd19217: duty=168; 15'd19218: duty=172; 15'd19219: duty=180; 15'd19220: duty=167; 15'd19221: duty=169; 15'd19222: duty=164; 15'd19223: duty=165;
15'd19224: duty=164; 15'd19225: duty=164; 15'd19226: duty=153; 15'd19227: duty=157; 15'd19228: duty=164; 15'd19229: duty=169; 15'd19230: duty=170; 15'd19231: duty=161;
15'd19232: duty=162; 15'd19233: duty=160; 15'd19234: duty=161; 15'd19235: duty=152; 15'd19236: duty=161; 15'd19237: duty=163; 15'd19238: duty=155; 15'd19239: duty=145;
15'd19240: duty=139; 15'd19241: duty=143; 15'd19242: duty=141; 15'd19243: duty=132; 15'd19244: duty=124; 15'd19245: duty=125; 15'd19246: duty=128; 15'd19247: duty=118;
15'd19248: duty=112; 15'd19249: duty=115; 15'd19250: duty=114; 15'd19251: duty=115; 15'd19252: duty=83; 15'd19253: duty=92; 15'd19254: duty=114; 15'd19255: duty=110;
15'd19256: duty=104; 15'd19257: duty=97; 15'd19258: duty=101; 15'd19259: duty=107; 15'd19260: duty=96; 15'd19261: duty=91; 15'd19262: duty=98; 15'd19263: duty=101;
15'd19264: duty=100; 15'd19265: duty=93; 15'd19266: duty=103; 15'd19267: duty=92; 15'd19268: duty=87; 15'd19269: duty=88; 15'd19270: duty=87; 15'd19271: duty=104;
15'd19272: duty=109; 15'd19273: duty=99; 15'd19274: duty=106; 15'd19275: duty=102; 15'd19276: duty=113; 15'd19277: duty=122; 15'd19278: duty=114; 15'd19279: duty=114;
15'd19280: duty=116; 15'd19281: duty=127; 15'd19282: duty=124; 15'd19283: duty=124; 15'd19284: duty=130; 15'd19285: duty=122; 15'd19286: duty=131; 15'd19287: duty=142;
15'd19288: duty=128; 15'd19289: duty=129; 15'd19290: duty=139; 15'd19291: duty=143; 15'd19292: duty=146; 15'd19293: duty=168; 15'd19294: duty=165; 15'd19295: duty=159;
15'd19296: duty=172; 15'd19297: duty=165; 15'd19298: duty=171; 15'd19299: duty=179; 15'd19300: duty=168; 15'd19301: duty=173; 15'd19302: duty=169; 15'd19303: duty=167;
15'd19304: duty=173; 15'd19305: duty=176; 15'd19306: duty=176; 15'd19307: duty=168; 15'd19308: duty=166; 15'd19309: duty=170; 15'd19310: duty=160; 15'd19311: duty=157;
15'd19312: duty=165; 15'd19313: duty=154; 15'd19314: duty=156; 15'd19315: duty=148; 15'd19316: duty=140; 15'd19317: duty=144; 15'd19318: duty=137; 15'd19319: duty=133;
15'd19320: duty=131; 15'd19321: duty=130; 15'd19322: duty=127; 15'd19323: duty=131; 15'd19324: duty=128; 15'd19325: duty=122; 15'd19326: duty=121; 15'd19327: duty=116;
15'd19328: duty=107; 15'd19329: duty=111; 15'd19330: duty=106; 15'd19331: duty=99; 15'd19332: duty=112; 15'd19333: duty=110; 15'd19334: duty=113; 15'd19335: duty=112;
15'd19336: duty=107; 15'd19337: duty=93; 15'd19338: duty=99; 15'd19339: duty=93; 15'd19340: duty=99; 15'd19341: duty=104; 15'd19342: duty=96; 15'd19343: duty=95;
15'd19344: duty=93; 15'd19345: duty=91; 15'd19346: duty=96; 15'd19347: duty=104; 15'd19348: duty=100; 15'd19349: duty=107; 15'd19350: duty=102; 15'd19351: duty=109;
15'd19352: duty=107; 15'd19353: duty=122; 15'd19354: duty=124; 15'd19355: duty=119; 15'd19356: duty=116; 15'd19357: duty=112; 15'd19358: duty=116; 15'd19359: duty=132;
15'd19360: duty=139; 15'd19361: duty=140; 15'd19362: duty=150; 15'd19363: duty=136; 15'd19364: duty=139; 15'd19365: duty=136; 15'd19366: duty=134; 15'd19367: duty=142;
15'd19368: duty=147; 15'd19369: duty=142; 15'd19370: duty=139; 15'd19371: duty=148; 15'd19372: duty=147; 15'd19373: duty=143; 15'd19374: duty=162; 15'd19375: duty=171;
15'd19376: duty=170; 15'd19377: duty=173; 15'd19378: duty=167; 15'd19379: duty=174; 15'd19380: duty=179; 15'd19381: duty=169; 15'd19382: duty=170; 15'd19383: duty=169;
15'd19384: duty=153; 15'd19385: duty=149; 15'd19386: duty=150; 15'd19387: duty=145; 15'd19388: duty=150; 15'd19389: duty=149; 15'd19390: duty=142; 15'd19391: duty=152;
15'd19392: duty=153; 15'd19393: duty=151; 15'd19394: duty=152; 15'd19395: duty=149; 15'd19396: duty=139; 15'd19397: duty=127; 15'd19398: duty=126; 15'd19399: duty=128;
15'd19400: duty=129; 15'd19401: duty=119; 15'd19402: duty=121; 15'd19403: duty=125; 15'd19404: duty=127; 15'd19405: duty=122; 15'd19406: duty=112; 15'd19407: duty=116;
15'd19408: duty=110; 15'd19409: duty=104; 15'd19410: duty=112; 15'd19411: duty=111; 15'd19412: duty=107; 15'd19413: duty=107; 15'd19414: duty=102; 15'd19415: duty=104;
15'd19416: duty=119; 15'd19417: duty=113; 15'd19418: duty=119; 15'd19419: duty=106; 15'd19420: duty=95; 15'd19421: duty=95; 15'd19422: duty=86; 15'd19423: duty=98;
15'd19424: duty=94; 15'd19425: duty=89; 15'd19426: duty=84; 15'd19427: duty=86; 15'd19428: duty=96; 15'd19429: duty=106; 15'd19430: duty=110; 15'd19431: duty=128;
15'd19432: duty=129; 15'd19433: duty=124; 15'd19434: duty=125; 15'd19435: duty=134; 15'd19436: duty=129; 15'd19437: duty=109; 15'd19438: duty=105; 15'd19439: duty=114;
15'd19440: duty=128; 15'd19441: duty=135; 15'd19442: duty=138; 15'd19443: duty=138; 15'd19444: duty=137; 15'd19445: duty=142; 15'd19446: duty=154; 15'd19447: duty=161;
15'd19448: duty=160; 15'd19449: duty=154; 15'd19450: duty=140; 15'd19451: duty=139; 15'd19452: duty=151; 15'd19453: duty=148; 15'd19454: duty=159; 15'd19455: duty=156;
15'd19456: duty=159; 15'd19457: duty=171; 15'd19458: duty=179; 15'd19459: duty=182; 15'd19460: duty=182; 15'd19461: duty=177; 15'd19462: duty=179; 15'd19463: duty=178;
15'd19464: duty=178; 15'd19465: duty=168; 15'd19466: duty=161; 15'd19467: duty=149; 15'd19468: duty=136; 15'd19469: duty=142; 15'd19470: duty=139; 15'd19471: duty=149;
15'd19472: duty=144; 15'd19473: duty=148; 15'd19474: duty=147; 15'd19475: duty=148; 15'd19476: duty=146; 15'd19477: duty=141; 15'd19478: duty=134; 15'd19479: duty=125;
15'd19480: duty=133; 15'd19481: duty=120; 15'd19482: duty=115; 15'd19483: duty=117; 15'd19484: duty=101; 15'd19485: duty=91; 15'd19486: duty=99; 15'd19487: duty=107;
15'd19488: duty=118; 15'd19489: duty=113; 15'd19490: duty=101; 15'd19491: duty=104; 15'd19492: duty=107; 15'd19493: duty=110; 15'd19494: duty=98; 15'd19495: duty=92;
15'd19496: duty=94; 15'd19497: duty=101; 15'd19498: duty=101; 15'd19499: duty=106; 15'd19500: duty=100; 15'd19501: duty=98; 15'd19502: duty=107; 15'd19503: duty=95;
15'd19504: duty=110; 15'd19505: duty=106; 15'd19506: duty=100; 15'd19507: duty=112; 15'd19508: duty=104; 15'd19509: duty=112; 15'd19510: duty=111; 15'd19511: duty=109;
15'd19512: duty=111; 15'd19513: duty=109; 15'd19514: duty=120; 15'd19515: duty=127; 15'd19516: duty=123; 15'd19517: duty=133; 15'd19518: duty=134; 15'd19519: duty=117;
15'd19520: duty=122; 15'd19521: duty=133; 15'd19522: duty=135; 15'd19523: duty=138; 15'd19524: duty=137; 15'd19525: duty=124; 15'd19526: duty=140; 15'd19527: duty=136;
15'd19528: duty=134; 15'd19529: duty=142; 15'd19530: duty=140; 15'd19531: duty=142; 15'd19532: duty=154; 15'd19533: duty=161; 15'd19534: duty=163; 15'd19535: duty=165;
15'd19536: duty=169; 15'd19537: duty=191; 15'd19538: duty=176; 15'd19539: duty=182; 15'd19540: duty=184; 15'd19541: duty=170; 15'd19542: duty=163; 15'd19543: duty=154;
15'd19544: duty=159; 15'd19545: duty=162; 15'd19546: duty=164; 15'd19547: duty=152; 15'd19548: duty=153; 15'd19549: duty=149; 15'd19550: duty=147; 15'd19551: duty=160;
15'd19552: duty=153; 15'd19553: duty=151; 15'd19554: duty=146; 15'd19555: duty=134; 15'd19556: duty=143; 15'd19557: duty=144; 15'd19558: duty=135; 15'd19559: duty=140;
15'd19560: duty=133; 15'd19561: duty=132; 15'd19562: duty=138; 15'd19563: duty=131; 15'd19564: duty=133; 15'd19565: duty=120; 15'd19566: duty=112; 15'd19567: duty=115;
15'd19568: duty=111; 15'd19569: duty=107; 15'd19570: duty=112; 15'd19571: duty=94; 15'd19572: duty=92; 15'd19573: duty=83; 15'd19574: duty=89; 15'd19575: duty=106;
15'd19576: duty=98; 15'd19577: duty=96; 15'd19578: duty=92; 15'd19579: duty=99; 15'd19580: duty=104; 15'd19581: duty=105; 15'd19582: duty=100; 15'd19583: duty=99;
15'd19584: duty=96; 15'd19585: duty=101; 15'd19586: duty=101; 15'd19587: duty=109; 15'd19588: duty=119; 15'd19589: duty=100; 15'd19590: duty=90; 15'd19591: duty=101;
15'd19592: duty=108; 15'd19593: duty=118; 15'd19594: duty=106; 15'd19595: duty=114; 15'd19596: duty=123; 15'd19597: duty=120; 15'd19598: duty=129; 15'd19599: duty=136;
15'd19600: duty=132; 15'd19601: duty=125; 15'd19602: duty=125; 15'd19603: duty=153; 15'd19604: duty=165; 15'd19605: duty=160; 15'd19606: duty=154; 15'd19607: duty=132;
15'd19608: duty=131; 15'd19609: duty=152; 15'd19610: duty=156; 15'd19611: duty=156; 15'd19612: duty=148; 15'd19613: duty=135; 15'd19614: duty=157; 15'd19615: duty=159;
15'd19616: duty=172; 15'd19617: duty=174; 15'd19618: duty=168; 15'd19619: duty=165; 15'd19620: duty=173; 15'd19621: duty=176; 15'd19622: duty=179; 15'd19623: duty=179;
15'd19624: duty=165; 15'd19625: duty=162; 15'd19626: duty=155; 15'd19627: duty=154; 15'd19628: duty=156; 15'd19629: duty=149; 15'd19630: duty=150; 15'd19631: duty=150;
15'd19632: duty=150; 15'd19633: duty=151; 15'd19634: duty=150; 15'd19635: duty=146; 15'd19636: duty=143; 15'd19637: duty=130; 15'd19638: duty=121; 15'd19639: duty=140;
15'd19640: duty=131; 15'd19641: duty=125; 15'd19642: duty=124; 15'd19643: duty=116; 15'd19644: duty=109; 15'd19645: duty=108; 15'd19646: duty=102; 15'd19647: duty=113;
15'd19648: duty=103; 15'd19649: duty=95; 15'd19650: duty=101; 15'd19651: duty=107; 15'd19652: duty=119; 15'd19653: duty=118; 15'd19654: duty=107; 15'd19655: duty=88;
15'd19656: duty=70; 15'd19657: duty=70; 15'd19658: duty=91; 15'd19659: duty=95; 15'd19660: duty=99; 15'd19661: duty=96; 15'd19662: duty=78; 15'd19663: duty=77;
15'd19664: duty=87; 15'd19665: duty=106; 15'd19666: duty=105; 15'd19667: duty=110; 15'd19668: duty=111; 15'd19669: duty=103; 15'd19670: duty=110; 15'd19671: duty=111;
15'd19672: duty=111; 15'd19673: duty=114; 15'd19674: duty=119; 15'd19675: duty=109; 15'd19676: duty=127; 15'd19677: duty=132; 15'd19678: duty=128; 15'd19679: duty=133;
15'd19680: duty=124; 15'd19681: duty=135; 15'd19682: duty=141; 15'd19683: duty=142; 15'd19684: duty=149; 15'd19685: duty=142; 15'd19686: duty=146; 15'd19687: duty=156;
15'd19688: duty=156; 15'd19689: duty=164; 15'd19690: duty=162; 15'd19691: duty=144; 15'd19692: duty=158; 15'd19693: duty=165; 15'd19694: duty=163; 15'd19695: duty=169;
15'd19696: duty=171; 15'd19697: duty=184; 15'd19698: duty=191; 15'd19699: duty=199; 15'd19700: duty=192; 15'd19701: duty=179; 15'd19702: duty=175; 15'd19703: duty=173;
15'd19704: duty=171; 15'd19705: duty=162; 15'd19706: duty=155; 15'd19707: duty=155; 15'd19708: duty=144; 15'd19709: duty=152; 15'd19710: duty=154; 15'd19711: duty=151;
15'd19712: duty=158; 15'd19713: duty=148; 15'd19714: duty=141; 15'd19715: duty=154; 15'd19716: duty=154; 15'd19717: duty=138; 15'd19718: duty=130; 15'd19719: duty=129;
15'd19720: duty=122; 15'd19721: duty=120; 15'd19722: duty=118; 15'd19723: duty=121; 15'd19724: duty=109; 15'd19725: duty=109; 15'd19726: duty=114; 15'd19727: duty=115;
15'd19728: duty=115; 15'd19729: duty=96; 15'd19730: duty=95; 15'd19731: duty=92; 15'd19732: duty=86; 15'd19733: duty=80; 15'd19734: duty=82; 15'd19735: duty=88;
15'd19736: duty=88; 15'd19737: duty=88; 15'd19738: duty=82; 15'd19739: duty=74; 15'd19740: duty=83; 15'd19741: duty=83; 15'd19742: duty=88; 15'd19743: duty=95;
15'd19744: duty=83; 15'd19745: duty=84; 15'd19746: duty=92; 15'd19747: duty=94; 15'd19748: duty=94; 15'd19749: duty=101; 15'd19750: duty=92; 15'd19751: duty=96;
15'd19752: duty=120; 15'd19753: duty=130; 15'd19754: duty=128; 15'd19755: duty=116; 15'd19756: duty=129; 15'd19757: duty=139; 15'd19758: duty=134; 15'd19759: duty=131;
15'd19760: duty=125; 15'd19761: duty=136; 15'd19762: duty=138; 15'd19763: duty=136; 15'd19764: duty=131; 15'd19765: duty=137; 15'd19766: duty=146; 15'd19767: duty=151;
15'd19768: duty=159; 15'd19769: duty=153; 15'd19770: duty=170; 15'd19771: duty=171; 15'd19772: duty=171; 15'd19773: duty=171; 15'd19774: duty=180; 15'd19775: duty=170;
15'd19776: duty=165; 15'd19777: duty=175; 15'd19778: duty=176; 15'd19779: duty=199; 15'd19780: duty=187; 15'd19781: duty=186; 15'd19782: duty=193; 15'd19783: duty=186;
15'd19784: duty=178; 15'd19785: duty=178; 15'd19786: duty=171; 15'd19787: duty=174; 15'd19788: duty=171; 15'd19789: duty=171; 15'd19790: duty=171; 15'd19791: duty=168;
15'd19792: duty=168; 15'd19793: duty=169; 15'd19794: duty=152; 15'd19795: duty=144; 15'd19796: duty=146; 15'd19797: duty=141; 15'd19798: duty=133; 15'd19799: duty=123;
15'd19800: duty=128; 15'd19801: duty=124; 15'd19802: duty=113; 15'd19803: duty=104; 15'd19804: duty=111; 15'd19805: duty=101; 15'd19806: duty=114; 15'd19807: duty=107;
15'd19808: duty=97; 15'd19809: duty=95; 15'd19810: duty=92; 15'd19811: duty=88; 15'd19812: duty=92; 15'd19813: duty=92; 15'd19814: duty=93; 15'd19815: duty=88;
15'd19816: duty=72; 15'd19817: duty=79; 15'd19818: duty=86; 15'd19819: duty=82; 15'd19820: duty=83; 15'd19821: duty=81; 15'd19822: duty=68; 15'd19823: duty=82;
15'd19824: duty=74; 15'd19825: duty=94; 15'd19826: duty=108; 15'd19827: duty=111; 15'd19828: duty=113; 15'd19829: duty=108; 15'd19830: duty=97; 15'd19831: duty=106;
15'd19832: duty=116; 15'd19833: duty=113; 15'd19834: duty=118; 15'd19835: duty=107; 15'd19836: duty=110; 15'd19837: duty=105; 15'd19838: duty=96; 15'd19839: duty=104;
15'd19840: duty=117; 15'd19841: duty=124; 15'd19842: duty=121; 15'd19843: duty=129; 15'd19844: duty=153; 15'd19845: duty=154; 15'd19846: duty=150; 15'd19847: duty=161;
15'd19848: duty=156; 15'd19849: duty=150; 15'd19850: duty=156; 15'd19851: duty=152; 15'd19852: duty=160; 15'd19853: duty=158; 15'd19854: duty=149; 15'd19855: duty=155;
15'd19856: duty=170; 15'd19857: duty=181; 15'd19858: duty=177; 15'd19859: duty=183; 15'd19860: duty=192; 15'd19861: duty=187; 15'd19862: duty=192; 15'd19863: duty=187;
15'd19864: duty=175; 15'd19865: duty=169; 15'd19866: duty=172; 15'd19867: duty=174; 15'd19868: duty=168; 15'd19869: duty=167; 15'd19870: duty=161; 15'd19871: duty=175;
15'd19872: duty=177; 15'd19873: duty=185; 15'd19874: duty=176; 15'd19875: duty=160; 15'd19876: duty=153; 15'd19877: duty=139; 15'd19878: duty=144; 15'd19879: duty=144;
15'd19880: duty=129; 15'd19881: duty=120; 15'd19882: duty=125; 15'd19883: duty=118; 15'd19884: duty=120; 15'd19885: duty=129; 15'd19886: duty=128; 15'd19887: duty=114;
15'd19888: duty=112; 15'd19889: duty=94; 15'd19890: duty=86; 15'd19891: duty=102; 15'd19892: duty=103; 15'd19893: duty=91; 15'd19894: duty=76; 15'd19895: duty=84;
15'd19896: duty=82; 15'd19897: duty=91; 15'd19898: duty=100; 15'd19899: duty=104; 15'd19900: duty=88; 15'd19901: duty=104; 15'd19902: duty=105; 15'd19903: duty=81;
15'd19904: duty=88; 15'd19905: duty=78; 15'd19906: duty=76; 15'd19907: duty=72; 15'd19908: duty=78; 15'd19909: duty=82; 15'd19910: duty=97; 15'd19911: duty=99;
15'd19912: duty=101; 15'd19913: duty=111; 15'd19914: duty=126; 15'd19915: duty=129; 15'd19916: duty=112; 15'd19917: duty=116; 15'd19918: duty=122; 15'd19919: duty=119;
15'd19920: duty=129; 15'd19921: duty=125; 15'd19922: duty=118; 15'd19923: duty=126; 15'd19924: duty=129; 15'd19925: duty=131; 15'd19926: duty=140; 15'd19927: duty=163;
15'd19928: duty=162; 15'd19929: duty=158; 15'd19930: duty=153; 15'd19931: duty=140; 15'd19932: duty=150; 15'd19933: duty=166; 15'd19934: duty=154; 15'd19935: duty=154;
15'd19936: duty=160; 15'd19937: duty=172; 15'd19938: duty=177; 15'd19939: duty=183; 15'd19940: duty=175; 15'd19941: duty=176; 15'd19942: duty=190; 15'd19943: duty=195;
15'd19944: duty=193; 15'd19945: duty=179; 15'd19946: duty=169; 15'd19947: duty=159; 15'd19948: duty=161; 15'd19949: duty=151; 15'd19950: duty=145; 15'd19951: duty=148;
15'd19952: duty=154; 15'd19953: duty=152; 15'd19954: duty=157; 15'd19955: duty=165; 15'd19956: duty=159; 15'd19957: duty=145; 15'd19958: duty=137; 15'd19959: duty=138;
15'd19960: duty=145; 15'd19961: duty=142; 15'd19962: duty=131; 15'd19963: duty=122; 15'd19964: duty=105; 15'd19965: duty=96; 15'd19966: duty=90; 15'd19967: duty=108;
15'd19968: duty=107; 15'd19969: duty=110; 15'd19970: duty=102; 15'd19971: duty=93; 15'd19972: duty=110; 15'd19973: duty=105; 15'd19974: duty=109; 15'd19975: duty=99;
15'd19976: duty=93; 15'd19977: duty=108; 15'd19978: duty=98; 15'd19979: duty=97; 15'd19980: duty=111; 15'd19981: duty=90; 15'd19982: duty=84; 15'd19983: duty=85;
15'd19984: duty=80; 15'd19985: duty=85; 15'd19986: duty=98; 15'd19987: duty=106; 15'd19988: duty=116; 15'd19989: duty=102; 15'd19990: duty=112; 15'd19991: duty=114;
15'd19992: duty=118; 15'd19993: duty=116; 15'd19994: duty=101; 15'd19995: duty=125; 15'd19996: duty=130; 15'd19997: duty=128; 15'd19998: duty=108; 15'd19999: duty=110;
15'd20000: duty=111; 15'd20001: duty=127; 15'd20002: duty=134; 15'd20003: duty=141; 15'd20004: duty=145; 15'd20005: duty=140; 15'd20006: duty=137; 15'd20007: duty=141;
15'd20008: duty=145; 15'd20009: duty=140; 15'd20010: duty=139; 15'd20011: duty=149; 15'd20012: duty=147; 15'd20013: duty=146; 15'd20014: duty=170; 15'd20015: duty=165;
15'd20016: duty=161; 15'd20017: duty=169; 15'd20018: duty=182; 15'd20019: duty=192; 15'd20020: duty=185; 15'd20021: duty=176; 15'd20022: duty=178; 15'd20023: duty=173;
15'd20024: duty=167; 15'd20025: duty=160; 15'd20026: duty=153; 15'd20027: duty=163; 15'd20028: duty=160; 15'd20029: duty=154; 15'd20030: duty=167; 15'd20031: duty=163;
15'd20032: duty=168; 15'd20033: duty=169; 15'd20034: duty=154; 15'd20035: duty=140; 15'd20036: duty=134; 15'd20037: duty=128; 15'd20038: duty=127; 15'd20039: duty=127;
15'd20040: duty=124; 15'd20041: duty=113; 15'd20042: duty=127; 15'd20043: duty=129; 15'd20044: duty=125; 15'd20045: duty=128; 15'd20046: duty=118; 15'd20047: duty=115;
15'd20048: duty=114; 15'd20049: duty=112; 15'd20050: duty=90; 15'd20051: duty=98; 15'd20052: duty=102; 15'd20053: duty=92; 15'd20054: duty=87; 15'd20055: duty=83;
15'd20056: duty=87; 15'd20057: duty=95; 15'd20058: duty=91; 15'd20059: duty=93; 15'd20060: duty=96; 15'd20061: duty=101; 15'd20062: duty=105; 15'd20063: duty=96;
15'd20064: duty=98; 15'd20065: duty=98; 15'd20066: duty=96; 15'd20067: duty=107; 15'd20068: duty=102; 15'd20069: duty=99; 15'd20070: duty=105; 15'd20071: duty=95;
15'd20072: duty=102; 15'd20073: duty=96; 15'd20074: duty=107; 15'd20075: duty=129; 15'd20076: duty=134; 15'd20077: duty=138; 15'd20078: duty=142; 15'd20079: duty=141;
15'd20080: duty=140; 15'd20081: duty=144; 15'd20082: duty=134; 15'd20083: duty=142; 15'd20084: duty=134; 15'd20085: duty=137; 15'd20086: duty=143; 15'd20087: duty=139;
15'd20088: duty=145; 15'd20089: duty=137; 15'd20090: duty=153; 15'd20091: duty=144; 15'd20092: duty=157; 15'd20093: duty=174; 15'd20094: duty=165; 15'd20095: duty=173;
15'd20096: duty=173; 15'd20097: duty=174; 15'd20098: duty=185; 15'd20099: duty=190; 15'd20100: duty=188; 15'd20101: duty=188; 15'd20102: duty=179; 15'd20103: duty=176;
15'd20104: duty=182; 15'd20105: duty=174; 15'd20106: duty=167; 15'd20107: duty=154; 15'd20108: duty=146; 15'd20109: duty=146; 15'd20110: duty=144; 15'd20111: duty=149;
15'd20112: duty=147; 15'd20113: duty=142; 15'd20114: duty=134; 15'd20115: duty=127; 15'd20116: duty=123; 15'd20117: duty=129; 15'd20118: duty=140; 15'd20119: duty=137;
15'd20120: duty=123; 15'd20121: duty=124; 15'd20122: duty=124; 15'd20123: duty=113; 15'd20124: duty=102; 15'd20125: duty=104; 15'd20126: duty=107; 15'd20127: duty=104;
15'd20128: duty=108; 15'd20129: duty=104; 15'd20130: duty=98; 15'd20131: duty=86; 15'd20132: duty=96; 15'd20133: duty=99; 15'd20134: duty=99; 15'd20135: duty=113;
15'd20136: duty=104; 15'd20137: duty=103; 15'd20138: duty=98; 15'd20139: duty=98; 15'd20140: duty=99; 15'd20141: duty=93; 15'd20142: duty=93; 15'd20143: duty=107;
15'd20144: duty=113; 15'd20145: duty=107; 15'd20146: duty=116; 15'd20147: duty=117; 15'd20148: duty=116; 15'd20149: duty=112; 15'd20150: duty=101; 15'd20151: duty=119;
15'd20152: duty=123; 15'd20153: duty=124; 15'd20154: duty=116; 15'd20155: duty=110; 15'd20156: duty=111; 15'd20157: duty=120; 15'd20158: duty=128; 15'd20159: duty=127;
15'd20160: duty=133; 15'd20161: duty=131; 15'd20162: duty=136; 15'd20163: duty=142; 15'd20164: duty=140; 15'd20165: duty=127; 15'd20166: duty=131; 15'd20167: duty=133;
15'd20168: duty=144; 15'd20169: duty=143; 15'd20170: duty=148; 15'd20171: duty=160; 15'd20172: duty=162; 15'd20173: duty=160; 15'd20174: duty=168; 15'd20175: duty=169;
15'd20176: duty=174; 15'd20177: duty=180; 15'd20178: duty=176; 15'd20179: duty=171; 15'd20180: duty=167; 15'd20181: duty=172; 15'd20182: duty=153; 15'd20183: duty=143;
15'd20184: duty=153; 15'd20185: duty=152; 15'd20186: duty=162; 15'd20187: duty=169; 15'd20188: duty=159; 15'd20189: duty=162; 15'd20190: duty=157; 15'd20191: duty=160;
15'd20192: duty=163; 15'd20193: duty=157; 15'd20194: duty=150; 15'd20195: duty=146; 15'd20196: duty=134; 15'd20197: duty=135; 15'd20198: duty=132; 15'd20199: duty=141;
15'd20200: duty=131; 15'd20201: duty=127; 15'd20202: duty=126; 15'd20203: duty=115; 15'd20204: duty=122; 15'd20205: duty=119; 15'd20206: duty=110; 15'd20207: duty=110;
15'd20208: duty=120; 15'd20209: duty=108; 15'd20210: duty=109; 15'd20211: duty=99; 15'd20212: duty=106; 15'd20213: duty=105; 15'd20214: duty=100; 15'd20215: duty=107;
15'd20216: duty=105; 15'd20217: duty=103; 15'd20218: duty=99; 15'd20219: duty=95; 15'd20220: duty=90; 15'd20221: duty=93; 15'd20222: duty=95; 15'd20223: duty=95;
15'd20224: duty=95; 15'd20225: duty=90; 15'd20226: duty=72; 15'd20227: duty=70; 15'd20228: duty=81; 15'd20229: duty=101; 15'd20230: duty=118; 15'd20231: duty=112;
15'd20232: duty=124; 15'd20233: duty=127; 15'd20234: duty=121; 15'd20235: duty=127; 15'd20236: duty=126; 15'd20237: duty=127; 15'd20238: duty=133; 15'd20239: duty=127;
15'd20240: duty=133; 15'd20241: duty=128; 15'd20242: duty=119; 15'd20243: duty=124; 15'd20244: duty=125; 15'd20245: duty=134; 15'd20246: duty=137; 15'd20247: duty=145;
15'd20248: duty=150; 15'd20249: duty=153; 15'd20250: duty=151; 15'd20251: duty=166; 15'd20252: duty=167; 15'd20253: duty=156; 15'd20254: duty=168; 15'd20255: duty=169;
15'd20256: duty=171; 15'd20257: duty=182; 15'd20258: duty=176; 15'd20259: duty=163; 15'd20260: duty=156; 15'd20261: duty=154; 15'd20262: duty=173; 15'd20263: duty=174;
15'd20264: duty=174; 15'd20265: duty=174; 15'd20266: duty=159; 15'd20267: duty=154; 15'd20268: duty=158; 15'd20269: duty=169; 15'd20270: duty=162; 15'd20271: duty=156;
15'd20272: duty=148; 15'd20273: duty=156; 15'd20274: duty=156; 15'd20275: duty=143; 15'd20276: duty=142; 15'd20277: duty=129; 15'd20278: duty=121; 15'd20279: duty=122;
15'd20280: duty=142; 15'd20281: duty=139; 15'd20282: duty=131; 15'd20283: duty=121; 15'd20284: duty=127; 15'd20285: duty=134; 15'd20286: duty=129; 15'd20287: duty=110;
15'd20288: duty=107; 15'd20289: duty=124; 15'd20290: duty=110; 15'd20291: duty=109; 15'd20292: duty=90; 15'd20293: duty=83; 15'd20294: duty=88; 15'd20295: duty=93;
15'd20296: duty=110; 15'd20297: duty=104; 15'd20298: duty=100; 15'd20299: duty=98; 15'd20300: duty=99; 15'd20301: duty=104; 15'd20302: duty=94; 15'd20303: duty=92;
15'd20304: duty=88; 15'd20305: duty=86; 15'd20306: duty=93; 15'd20307: duty=101; 15'd20308: duty=99; 15'd20309: duty=92; 15'd20310: duty=96; 15'd20311: duty=99;
15'd20312: duty=103; 15'd20313: duty=106; 15'd20314: duty=113; 15'd20315: duty=115; 15'd20316: duty=116; 15'd20317: duty=107; 15'd20318: duty=110; 15'd20319: duty=117;
15'd20320: duty=113; 15'd20321: duty=121; 15'd20322: duty=128; 15'd20323: duty=126; 15'd20324: duty=132; 15'd20325: duty=130; 15'd20326: duty=133; 15'd20327: duty=145;
15'd20328: duty=150; 15'd20329: duty=148; 15'd20330: duty=148; 15'd20331: duty=158; 15'd20332: duty=169; 15'd20333: duty=173; 15'd20334: duty=176; 15'd20335: duty=183;
15'd20336: duty=184; 15'd20337: duty=184; 15'd20338: duty=177; 15'd20339: duty=173; 15'd20340: duty=168; 15'd20341: duty=170; 15'd20342: duty=172; 15'd20343: duty=167;
15'd20344: duty=163; 15'd20345: duty=162; 15'd20346: duty=163; 15'd20347: duty=162; 15'd20348: duty=160; 15'd20349: duty=157; 15'd20350: duty=162; 15'd20351: duty=164;
15'd20352: duty=157; 15'd20353: duty=157; 15'd20354: duty=156; 15'd20355: duty=148; 15'd20356: duty=145; 15'd20357: duty=145; 15'd20358: duty=143; 15'd20359: duty=134;
15'd20360: duty=135; 15'd20361: duty=141; 15'd20362: duty=144; 15'd20363: duty=139; 15'd20364: duty=120; 15'd20365: duty=131; 15'd20366: duty=126; 15'd20367: duty=118;
15'd20368: duty=119; 15'd20369: duty=109; 15'd20370: duty=109; 15'd20371: duty=107; 15'd20372: duty=110; 15'd20373: duty=103; 15'd20374: duty=90; 15'd20375: duty=86;
15'd20376: duty=93; 15'd20377: duty=95; 15'd20378: duty=99; 15'd20379: duty=101; 15'd20380: duty=92; 15'd20381: duty=92; 15'd20382: duty=91; 15'd20383: duty=90;
15'd20384: duty=96; 15'd20385: duty=95; 15'd20386: duty=85; 15'd20387: duty=84; 15'd20388: duty=84; 15'd20389: duty=82; 15'd20390: duty=95; 15'd20391: duty=98;
15'd20392: duty=105; 15'd20393: duty=113; 15'd20394: duty=115; 15'd20395: duty=116; 15'd20396: duty=112; 15'd20397: duty=124; 15'd20398: duty=115; 15'd20399: duty=118;
15'd20400: duty=122; 15'd20401: duty=121; 15'd20402: duty=130; 15'd20403: duty=125; 15'd20404: duty=136; 15'd20405: duty=139; 15'd20406: duty=137; 15'd20407: duty=142;
15'd20408: duty=147; 15'd20409: duty=150; 15'd20410: duty=150; 15'd20411: duty=148; 15'd20412: duty=151; 15'd20413: duty=161; 15'd20414: duty=162; 15'd20415: duty=165;
15'd20416: duty=166; 15'd20417: duty=171; 15'd20418: duty=171; 15'd20419: duty=171; 15'd20420: duty=171; 15'd20421: duty=173; 15'd20422: duty=159; 15'd20423: duty=156;
15'd20424: duty=160; 15'd20425: duty=148; 15'd20426: duty=154; 15'd20427: duty=156; 15'd20428: duty=151; 15'd20429: duty=153; 15'd20430: duty=157; 15'd20431: duty=171;
15'd20432: duty=168; 15'd20433: duty=158; 15'd20434: duty=160; 15'd20435: duty=154; 15'd20436: duty=142; 15'd20437: duty=145; 15'd20438: duty=142; 15'd20439: duty=139;
15'd20440: duty=136; 15'd20441: duty=128; 15'd20442: duty=131; 15'd20443: duty=125; 15'd20444: duty=124; 15'd20445: duty=121; 15'd20446: duty=121; 15'd20447: duty=118;
15'd20448: duty=117; 15'd20449: duty=110; 15'd20450: duty=125; 15'd20451: duty=116; 15'd20452: duty=113; 15'd20453: duty=117; 15'd20454: duty=107; 15'd20455: duty=108;
15'd20456: duty=105; 15'd20457: duty=108; 15'd20458: duty=102; 15'd20459: duty=96; 15'd20460: duty=102; 15'd20461: duty=106; 15'd20462: duty=109; 15'd20463: duty=107;
15'd20464: duty=115; 15'd20465: duty=115; 15'd20466: duty=115; 15'd20467: duty=107; 15'd20468: duty=105; 15'd20469: duty=90; 15'd20470: duty=91; 15'd20471: duty=95;
15'd20472: duty=88; 15'd20473: duty=104; 15'd20474: duty=108; 15'd20475: duty=113; 15'd20476: duty=116; 15'd20477: duty=118; 15'd20478: duty=115; 15'd20479: duty=128;
15'd20480: duty=119; 15'd20481: duty=134; 15'd20482: duty=135; 15'd20483: duty=131; 15'd20484: duty=137; 15'd20485: duty=130; 15'd20486: duty=130; 15'd20487: duty=133;
15'd20488: duty=131; 15'd20489: duty=136; 15'd20490: duty=146; 15'd20491: duty=150; 15'd20492: duty=156; 15'd20493: duty=157; 15'd20494: duty=166; 15'd20495: duty=167;
15'd20496: duty=176; 15'd20497: duty=170; 15'd20498: duty=151; 15'd20499: duty=142; 15'd20500: duty=154; 15'd20501: duty=165; 15'd20502: duty=166; 15'd20503: duty=157;
15'd20504: duty=160; 15'd20505: duty=153; 15'd20506: duty=154; 15'd20507: duty=170; 15'd20508: duty=171; 15'd20509: duty=167; 15'd20510: duty=154; 15'd20511: duty=145;
15'd20512: duty=141; 15'd20513: duty=144; 15'd20514: duty=139; 15'd20515: duty=137; 15'd20516: duty=134; 15'd20517: duty=139; 15'd20518: duty=150; 15'd20519: duty=148;
15'd20520: duty=143; 15'd20521: duty=136; 15'd20522: duty=131; 15'd20523: duty=122; 15'd20524: duty=113; 15'd20525: duty=116; 15'd20526: duty=121; 15'd20527: duty=115;
15'd20528: duty=94; 15'd20529: duty=93; 15'd20530: duty=101; 15'd20531: duty=102; 15'd20532: duty=105; 15'd20533: duty=104; 15'd20534: duty=116; 15'd20535: duty=112;
15'd20536: duty=104; 15'd20537: duty=102; 15'd20538: duty=110; 15'd20539: duty=104; 15'd20540: duty=110; 15'd20541: duty=107; 15'd20542: duty=105; 15'd20543: duty=112;
15'd20544: duty=102; 15'd20545: duty=107; 15'd20546: duty=101; 15'd20547: duty=98; 15'd20548: duty=107; 15'd20549: duty=106; 15'd20550: duty=110; 15'd20551: duty=124;
15'd20552: duty=108; 15'd20553: duty=115; 15'd20554: duty=114; 15'd20555: duty=118; 15'd20556: duty=124; 15'd20557: duty=121; 15'd20558: duty=118; 15'd20559: duty=134;
15'd20560: duty=136; 15'd20561: duty=121; 15'd20562: duty=128; 15'd20563: duty=128; 15'd20564: duty=134; 15'd20565: duty=142; 15'd20566: duty=159; 15'd20567: duty=156;
15'd20568: duty=162; 15'd20569: duty=155; 15'd20570: duty=159; 15'd20571: duty=160; 15'd20572: duty=160; 15'd20573: duty=162; 15'd20574: duty=162; 15'd20575: duty=162;
15'd20576: duty=165; 15'd20577: duty=169; 15'd20578: duty=173; 15'd20579: duty=171; 15'd20580: duty=164; 15'd20581: duty=162; 15'd20582: duty=158; 15'd20583: duty=168;
15'd20584: duty=169; 15'd20585: duty=164; 15'd20586: duty=159; 15'd20587: duty=154; 15'd20588: duty=147; 15'd20589: duty=146; 15'd20590: duty=149; 15'd20591: duty=147;
15'd20592: duty=138; 15'd20593: duty=138; 15'd20594: duty=135; 15'd20595: duty=134; 15'd20596: duty=127; 15'd20597: duty=130; 15'd20598: duty=127; 15'd20599: duty=123;
15'd20600: duty=120; 15'd20601: duty=123; 15'd20602: duty=120; 15'd20603: duty=114; 15'd20604: duty=117; 15'd20605: duty=111; 15'd20606: duty=114; 15'd20607: duty=102;
15'd20608: duty=100; 15'd20609: duty=103; 15'd20610: duty=103; 15'd20611: duty=104; 15'd20612: duty=98; 15'd20613: duty=97; 15'd20614: duty=102; 15'd20615: duty=97;
15'd20616: duty=92; 15'd20617: duty=77; 15'd20618: duty=72; 15'd20619: duty=79; 15'd20620: duty=90; 15'd20621: duty=99; 15'd20622: duty=105; 15'd20623: duty=101;
15'd20624: duty=107; 15'd20625: duty=111; 15'd20626: duty=112; 15'd20627: duty=116; 15'd20628: duty=115; 15'd20629: duty=111; 15'd20630: duty=107; 15'd20631: duty=113;
15'd20632: duty=112; 15'd20633: duty=119; 15'd20634: duty=115; 15'd20635: duty=121; 15'd20636: duty=122; 15'd20637: duty=129; 15'd20638: duty=143; 15'd20639: duty=145;
15'd20640: duty=139; 15'd20641: duty=134; 15'd20642: duty=136; 15'd20643: duty=148; 15'd20644: duty=156; 15'd20645: duty=159; 15'd20646: duty=160; 15'd20647: duty=162;
15'd20648: duty=176; 15'd20649: duty=185; 15'd20650: duty=190; 15'd20651: duty=193; 15'd20652: duty=189; 15'd20653: duty=181; 15'd20654: duty=173; 15'd20655: duty=167;
15'd20656: duty=171; 15'd20657: duty=165; 15'd20658: duty=154; 15'd20659: duty=148; 15'd20660: duty=154; 15'd20661: duty=164; 15'd20662: duty=169; 15'd20663: duty=161;
15'd20664: duty=152; 15'd20665: duty=156; 15'd20666: duty=162; 15'd20667: duty=162; 15'd20668: duty=160; 15'd20669: duty=163; 15'd20670: duty=149; 15'd20671: duty=142;
15'd20672: duty=140; 15'd20673: duty=132; 15'd20674: duty=137; 15'd20675: duty=127; 15'd20676: duty=122; 15'd20677: duty=122; 15'd20678: duty=125; 15'd20679: duty=133;
15'd20680: duty=122; 15'd20681: duty=120; 15'd20682: duty=115; 15'd20683: duty=101; 15'd20684: duty=97; 15'd20685: duty=85; 15'd20686: duty=93; 15'd20687: duty=106;
15'd20688: duty=94; 15'd20689: duty=78; 15'd20690: duty=91; 15'd20691: duty=91; 15'd20692: duty=85; 15'd20693: duty=91; 15'd20694: duty=80; 15'd20695: duty=88;
15'd20696: duty=93; 15'd20697: duty=104; 15'd20698: duty=110; 15'd20699: duty=100; 15'd20700: duty=97; 15'd20701: duty=87; 15'd20702: duty=82; 15'd20703: duty=106;
15'd20704: duty=116; 15'd20705: duty=102; 15'd20706: duty=95; 15'd20707: duty=95; 15'd20708: duty=99; 15'd20709: duty=110; 15'd20710: duty=110; 15'd20711: duty=117;
15'd20712: duty=131; 15'd20713: duty=131; 15'd20714: duty=141; 15'd20715: duty=137; 15'd20716: duty=129; 15'd20717: duty=131; 15'd20718: duty=133; 15'd20719: duty=137;
15'd20720: duty=139; 15'd20721: duty=152; 15'd20722: duty=157; 15'd20723: duty=149; 15'd20724: duty=151; 15'd20725: duty=154; 15'd20726: duty=158; 15'd20727: duty=172;
15'd20728: duty=161; 15'd20729: duty=161; 15'd20730: duty=176; 15'd20731: duty=176; 15'd20732: duty=179; 15'd20733: duty=174; 15'd20734: duty=168; 15'd20735: duty=176;
15'd20736: duty=183; 15'd20737: duty=180; 15'd20738: duty=179; 15'd20739: duty=169; 15'd20740: duty=168; 15'd20741: duty=171; 15'd20742: duty=165; 15'd20743: duty=162;
15'd20744: duty=159; 15'd20745: duty=144; 15'd20746: duty=148; 15'd20747: duty=150; 15'd20748: duty=143; 15'd20749: duty=144; 15'd20750: duty=143; 15'd20751: duty=130;
15'd20752: duty=125; 15'd20753: duty=131; 15'd20754: duty=124; 15'd20755: duty=123; 15'd20756: duty=122; 15'd20757: duty=118; 15'd20758: duty=122; 15'd20759: duty=121;
15'd20760: duty=117; 15'd20761: duty=113; 15'd20762: duty=99; 15'd20763: duty=100; 15'd20764: duty=93; 15'd20765: duty=90; 15'd20766: duty=104; 15'd20767: duty=109;
15'd20768: duty=101; 15'd20769: duty=92; 15'd20770: duty=88; 15'd20771: duty=86; 15'd20772: duty=93; 15'd20773: duty=96; 15'd20774: duty=98; 15'd20775: duty=100;
15'd20776: duty=105; 15'd20777: duty=113; 15'd20778: duty=102; 15'd20779: duty=115; 15'd20780: duty=121; 15'd20781: duty=102; 15'd20782: duty=96; 15'd20783: duty=91;
15'd20784: duty=92; 15'd20785: duty=108; 15'd20786: duty=124; 15'd20787: duty=117; 15'd20788: duty=116; 15'd20789: duty=121; 15'd20790: duty=125; 15'd20791: duty=129;
15'd20792: duty=126; 15'd20793: duty=122; 15'd20794: duty=128; 15'd20795: duty=129; 15'd20796: duty=131; 15'd20797: duty=136; 15'd20798: duty=139; 15'd20799: duty=136;
15'd20800: duty=133; 15'd20801: duty=136; 15'd20802: duty=149; 15'd20803: duty=153; 15'd20804: duty=150; 15'd20805: duty=165; 15'd20806: duty=168; 15'd20807: duty=177;
15'd20808: duty=174; 15'd20809: duty=168; 15'd20810: duty=176; 15'd20811: duty=168; 15'd20812: duty=174; 15'd20813: duty=168; 15'd20814: duty=160; 15'd20815: duty=154;
15'd20816: duty=152; 15'd20817: duty=153; 15'd20818: duty=163; 15'd20819: duty=165; 15'd20820: duty=162; 15'd20821: duty=171; 15'd20822: duty=157; 15'd20823: duty=168;
15'd20824: duty=170; 15'd20825: duty=170; 15'd20826: duty=168; 15'd20827: duty=158; 15'd20828: duty=146; 15'd20829: duty=144; 15'd20830: duty=145; 15'd20831: duty=134;
15'd20832: duty=135; 15'd20833: duty=117; 15'd20834: duty=111; 15'd20835: duty=109; 15'd20836: duty=119; 15'd20837: duty=115; 15'd20838: duty=120; 15'd20839: duty=104;
15'd20840: duty=111; 15'd20841: duty=128; 15'd20842: duty=111; 15'd20843: duty=108; 15'd20844: duty=86; 15'd20845: duty=93; 15'd20846: duty=94; 15'd20847: duty=92;
15'd20848: duty=83; 15'd20849: duty=83; 15'd20850: duty=77; 15'd20851: duty=80; 15'd20852: duty=102; 15'd20853: duty=98; 15'd20854: duty=108; 15'd20855: duty=104;
15'd20856: duty=96; 15'd20857: duty=84; 15'd20858: duty=79; 15'd20859: duty=78; 15'd20860: duty=87; 15'd20861: duty=107; 15'd20862: duty=114; 15'd20863: duty=127;
15'd20864: duty=124; 15'd20865: duty=116; 15'd20866: duty=118; 15'd20867: duty=125; 15'd20868: duty=127; 15'd20869: duty=126; 15'd20870: duty=134; 15'd20871: duty=133;
15'd20872: duty=130; 15'd20873: duty=130; 15'd20874: duty=136; 15'd20875: duty=139; 15'd20876: duty=134; 15'd20877: duty=137; 15'd20878: duty=139; 15'd20879: duty=146;
15'd20880: duty=164; 15'd20881: duty=157; 15'd20882: duty=156; 15'd20883: duty=153; 15'd20884: duty=156; 15'd20885: duty=166; 15'd20886: duty=167; 15'd20887: duty=168;
15'd20888: duty=171; 15'd20889: duty=172; 15'd20890: duty=167; 15'd20891: duty=175; 15'd20892: duty=176; 15'd20893: duty=176; 15'd20894: duty=168; 15'd20895: duty=171;
15'd20896: duty=171; 15'd20897: duty=169; 15'd20898: duty=167; 15'd20899: duty=159; 15'd20900: duty=158; 15'd20901: duty=159; 15'd20902: duty=158; 15'd20903: duty=148;
15'd20904: duty=156; 15'd20905: duty=155; 15'd20906: duty=136; 15'd20907: duty=145; 15'd20908: duty=142; 15'd20909: duty=138; 15'd20910: duty=143; 15'd20911: duty=132;
15'd20912: duty=128; 15'd20913: duty=119; 15'd20914: duty=124; 15'd20915: duty=124; 15'd20916: duty=118; 15'd20917: duty=111; 15'd20918: duty=98; 15'd20919: duty=99;
15'd20920: duty=101; 15'd20921: duty=95; 15'd20922: duty=96; 15'd20923: duty=96; 15'd20924: duty=95; 15'd20925: duty=94; 15'd20926: duty=103; 15'd20927: duty=102;
15'd20928: duty=83; 15'd20929: duty=79; 15'd20930: duty=87; 15'd20931: duty=101; 15'd20932: duty=98; 15'd20933: duty=90; 15'd20934: duty=89; 15'd20935: duty=96;
15'd20936: duty=101; 15'd20937: duty=99; 15'd20938: duty=99; 15'd20939: duty=99; 15'd20940: duty=104; 15'd20941: duty=104; 15'd20942: duty=104; 15'd20943: duty=115;
15'd20944: duty=113; 15'd20945: duty=115; 15'd20946: duty=108; 15'd20947: duty=115; 15'd20948: duty=126; 15'd20949: duty=127; 15'd20950: duty=127; 15'd20951: duty=128;
15'd20952: duty=143; 15'd20953: duty=130; 15'd20954: duty=139; 15'd20955: duty=137; 15'd20956: duty=145; 15'd20957: duty=148; 15'd20958: duty=149; 15'd20959: duty=161;
15'd20960: duty=153; 15'd20961: duty=156; 15'd20962: duty=148; 15'd20963: duty=151; 15'd20964: duty=163; 15'd20965: duty=177; 15'd20966: duty=183; 15'd20967: duty=191;
15'd20968: duty=183; 15'd20969: duty=179; 15'd20970: duty=177; 15'd20971: duty=172; 15'd20972: duty=177; 15'd20973: duty=167; 15'd20974: duty=169; 15'd20975: duty=168;
15'd20976: duty=169; 15'd20977: duty=171; 15'd20978: duty=165; 15'd20979: duty=150; 15'd20980: duty=140; 15'd20981: duty=142; 15'd20982: duty=148; 15'd20983: duty=154;
15'd20984: duty=154; 15'd20985: duty=154; 15'd20986: duty=148; 15'd20987: duty=140; 15'd20988: duty=140; 15'd20989: duty=145; 15'd20990: duty=135; 15'd20991: duty=128;
15'd20992: duty=129; 15'd20993: duty=128; 15'd20994: duty=130; 15'd20995: duty=121; 15'd20996: duty=111; 15'd20997: duty=102; 15'd20998: duty=90; 15'd20999: duty=102;
15'd21000: duty=105; 15'd21001: duty=110; 15'd21002: duty=109; 15'd21003: duty=101; 15'd21004: duty=93; 15'd21005: duty=79; 15'd21006: duty=90; 15'd21007: duty=96;
15'd21008: duty=101; 15'd21009: duty=96; 15'd21010: duty=93; 15'd21011: duty=92; 15'd21012: duty=88; 15'd21013: duty=89; 15'd21014: duty=81; 15'd21015: duty=79;
15'd21016: duty=82; 15'd21017: duty=96; 15'd21018: duty=97; 15'd21019: duty=96; 15'd21020: duty=98; 15'd21021: duty=93; 15'd21022: duty=94; 15'd21023: duty=106;
15'd21024: duty=110; 15'd21025: duty=110; 15'd21026: duty=110; 15'd21027: duty=115; 15'd21028: duty=128; 15'd21029: duty=124; 15'd21030: duty=123; 15'd21031: duty=136;
15'd21032: duty=139; 15'd21033: duty=148; 15'd21034: duty=155; 15'd21035: duty=144; 15'd21036: duty=137; 15'd21037: duty=139; 15'd21038: duty=143; 15'd21039: duty=144;
15'd21040: duty=149; 15'd21041: duty=150; 15'd21042: duty=160; 15'd21043: duty=162; 15'd21044: duty=166; 15'd21045: duty=179; 15'd21046: duty=182; 15'd21047: duty=182;
15'd21048: duty=188; 15'd21049: duty=184; 15'd21050: duty=180; 15'd21051: duty=187; 15'd21052: duty=180; 15'd21053: duty=182; 15'd21054: duty=173; 15'd21055: duty=159;
15'd21056: duty=163; 15'd21057: duty=159; 15'd21058: duty=162; 15'd21059: duty=169; 15'd21060: duty=170; 15'd21061: duty=165; 15'd21062: duty=168; 15'd21063: duty=168;
15'd21064: duty=167; 15'd21065: duty=154; 15'd21066: duty=150; 15'd21067: duty=149; 15'd21068: duty=130; 15'd21069: duty=136; 15'd21070: duty=130; 15'd21071: duty=131;
15'd21072: duty=130; 15'd21073: duty=125; 15'd21074: duty=119; 15'd21075: duty=108; 15'd21076: duty=112; 15'd21077: duty=108; 15'd21078: duty=101; 15'd21079: duty=90;
15'd21080: duty=100; 15'd21081: duty=100; 15'd21082: duty=92; 15'd21083: duty=100; 15'd21084: duty=100; 15'd21085: duty=96; 15'd21086: duty=103; 15'd21087: duty=98;
15'd21088: duty=98; 15'd21089: duty=97; 15'd21090: duty=87; 15'd21091: duty=78; 15'd21092: duty=84; 15'd21093: duty=99; 15'd21094: duty=104; 15'd21095: duty=92;
15'd21096: duty=99; 15'd21097: duty=101; 15'd21098: duty=101; 15'd21099: duty=105; 15'd21100: duty=100; 15'd21101: duty=101; 15'd21102: duty=104; 15'd21103: duty=104;
15'd21104: duty=95; 15'd21105: duty=98; 15'd21106: duty=85; 15'd21107: duty=101; 15'd21108: duty=108; 15'd21109: duty=110; 15'd21110: duty=113; 15'd21111: duty=128;
15'd21112: duty=146; 15'd21113: duty=139; 15'd21114: duty=146; 15'd21115: duty=144; 15'd21116: duty=144; 15'd21117: duty=141; 15'd21118: duty=147; 15'd21119: duty=148;
15'd21120: duty=152; 15'd21121: duty=151; 15'd21122: duty=153; 15'd21123: duty=164; 15'd21124: duty=170; 15'd21125: duty=173; 15'd21126: duty=182; 15'd21127: duty=177;
15'd21128: duty=176; 15'd21129: duty=181; 15'd21130: duty=167; 15'd21131: duty=167; 15'd21132: duty=165; 15'd21133: duty=167; 15'd21134: duty=168; 15'd21135: duty=171;
15'd21136: duty=167; 15'd21137: duty=171; 15'd21138: duty=177; 15'd21139: duty=168; 15'd21140: duty=163; 15'd21141: duty=170; 15'd21142: duty=161; 15'd21143: duty=151;
15'd21144: duty=157; 15'd21145: duty=152; 15'd21146: duty=153; 15'd21147: duty=148; 15'd21148: duty=148; 15'd21149: duty=145; 15'd21150: duty=134; 15'd21151: duty=140;
15'd21152: duty=131; 15'd21153: duty=125; 15'd21154: duty=136; 15'd21155: duty=122; 15'd21156: duty=115; 15'd21157: duty=110; 15'd21158: duty=104; 15'd21159: duty=102;
15'd21160: duty=100; 15'd21161: duty=94; 15'd21162: duty=90; 15'd21163: duty=83; 15'd21164: duty=83; 15'd21165: duty=94; 15'd21166: duty=84; 15'd21167: duty=85;
15'd21168: duty=98; 15'd21169: duty=94; 15'd21170: duty=95; 15'd21171: duty=99; 15'd21172: duty=87; 15'd21173: duty=104; 15'd21174: duty=95; 15'd21175: duty=76;
15'd21176: duty=81; 15'd21177: duty=76; 15'd21178: duty=89; 15'd21179: duty=99; 15'd21180: duty=98; 15'd21181: duty=102; 15'd21182: duty=115; 15'd21183: duty=106;
15'd21184: duty=110; 15'd21185: duty=110; 15'd21186: duty=110; 15'd21187: duty=128; 15'd21188: duty=133; 15'd21189: duty=134; 15'd21190: duty=140; 15'd21191: duty=134;
15'd21192: duty=123; 15'd21193: duty=126; 15'd21194: duty=128; 15'd21195: duty=148; 15'd21196: duty=148; 15'd21197: duty=136; 15'd21198: duty=133; 15'd21199: duty=142;
15'd21200: duty=163; 15'd21201: duty=165; 15'd21202: duty=163; 15'd21203: duty=162; 15'd21204: duty=168; 15'd21205: duty=170; 15'd21206: duty=182; 15'd21207: duty=192;
15'd21208: duty=187; 15'd21209: duty=185; 15'd21210: duty=177; 15'd21211: duty=166; 15'd21212: duty=164; 15'd21213: duty=163; 15'd21214: duty=162; 15'd21215: duty=164;
15'd21216: duty=161; 15'd21217: duty=166; 15'd21218: duty=162; 15'd21219: duty=165; 15'd21220: duty=163; 15'd21221: duty=161; 15'd21222: duty=162; 15'd21223: duty=161;
15'd21224: duty=167; 15'd21225: duty=161; 15'd21226: duty=155; 15'd21227: duty=146; 15'd21228: duty=139; 15'd21229: duty=136; 15'd21230: duty=130; 15'd21231: duty=122;
15'd21232: duty=117; 15'd21233: duty=123; 15'd21234: duty=122; 15'd21235: duty=114; 15'd21236: duty=106; 15'd21237: duty=109; 15'd21238: duty=111; 15'd21239: duty=106;
15'd21240: duty=114; 15'd21241: duty=108; 15'd21242: duty=97; 15'd21243: duty=102; 15'd21244: duty=95; 15'd21245: duty=103; 15'd21246: duty=103; 15'd21247: duty=80;
15'd21248: duty=83; 15'd21249: duty=83; 15'd21250: duty=81; 15'd21251: duty=91; 15'd21252: duty=95; 15'd21253: duty=103; 15'd21254: duty=103; 15'd21255: duty=96;
15'd21256: duty=97; 15'd21257: duty=96; 15'd21258: duty=100; 15'd21259: duty=108; 15'd21260: duty=100; 15'd21261: duty=98; 15'd21262: duty=97; 15'd21263: duty=93;
15'd21264: duty=120; 15'd21265: duty=119; 15'd21266: duty=121; 15'd21267: duty=124; 15'd21268: duty=117; 15'd21269: duty=125; 15'd21270: duty=130; 15'd21271: duty=130;
15'd21272: duty=126; 15'd21273: duty=115; 15'd21274: duty=121; 15'd21275: duty=126; 15'd21276: duty=128; 15'd21277: duty=147; 15'd21278: duty=148; 15'd21279: duty=149;
15'd21280: duty=166; 15'd21281: duty=174; 15'd21282: duty=166; 15'd21283: duty=181; 15'd21284: duty=180; 15'd21285: duty=179; 15'd21286: duty=180; 15'd21287: duty=179;
15'd21288: duty=171; 15'd21289: duty=164; 15'd21290: duty=163; 15'd21291: duty=167; 15'd21292: duty=170; 15'd21293: duty=171; 15'd21294: duty=176; 15'd21295: duty=162;
15'd21296: duty=163; 15'd21297: duty=171; 15'd21298: duty=163; 15'd21299: duty=161; 15'd21300: duty=159; 15'd21301: duty=155; 15'd21302: duty=144; 15'd21303: duty=144;
15'd21304: duty=136; 15'd21305: duty=139; 15'd21306: duty=143; 15'd21307: duty=127; 15'd21308: duty=128; 15'd21309: duty=114; 15'd21310: duty=125; 15'd21311: duty=135;
15'd21312: duty=126; 15'd21313: duty=123; 15'd21314: duty=123; 15'd21315: duty=115; 15'd21316: duty=111; 15'd21317: duty=108; 15'd21318: duty=115; 15'd21319: duty=114;
15'd21320: duty=105; 15'd21321: duty=103; 15'd21322: duty=102; 15'd21323: duty=94; 15'd21324: duty=85; 15'd21325: duty=82; 15'd21326: duty=82; 15'd21327: duty=86;
15'd21328: duty=85; 15'd21329: duty=88; 15'd21330: duty=91; 15'd21331: duty=86; 15'd21332: duty=100; 15'd21333: duty=113; 15'd21334: duty=113; 15'd21335: duty=111;
15'd21336: duty=101; 15'd21337: duty=103; 15'd21338: duty=113; 15'd21339: duty=124; 15'd21340: duty=127; 15'd21341: duty=113; 15'd21342: duty=93; 15'd21343: duty=104;
15'd21344: duty=116; 15'd21345: duty=127; 15'd21346: duty=127; 15'd21347: duty=128; 15'd21348: duty=126; 15'd21349: duty=131; 15'd21350: duty=122; 15'd21351: duty=134;
15'd21352: duty=133; 15'd21353: duty=135; 15'd21354: duty=143; 15'd21355: duty=148; 15'd21356: duty=157; 15'd21357: duty=154; 15'd21358: duty=165; 15'd21359: duty=170;
15'd21360: duty=173; 15'd21361: duty=164; 15'd21362: duty=175; 15'd21363: duty=175; 15'd21364: duty=164; 15'd21365: duty=166; 15'd21366: duty=173; 15'd21367: duty=172;
15'd21368: duty=170; 15'd21369: duty=162; 15'd21370: duty=161; 15'd21371: duty=167; 15'd21372: duty=165; 15'd21373: duty=163; 15'd21374: duty=165; 15'd21375: duty=164;
15'd21376: duty=161; 15'd21377: duty=161; 15'd21378: duty=150; 15'd21379: duty=152; 15'd21380: duty=147; 15'd21381: duty=137; 15'd21382: duty=139; 15'd21383: duty=127;
15'd21384: duty=127; 15'd21385: duty=124; 15'd21386: duty=124; 15'd21387: duty=126; 15'd21388: duty=129; 15'd21389: duty=125; 15'd21390: duty=124; 15'd21391: duty=118;
15'd21392: duty=114; 15'd21393: duty=113; 15'd21394: duty=111; 15'd21395: duty=118; 15'd21396: duty=112; 15'd21397: duty=112; 15'd21398: duty=97; 15'd21399: duty=93;
15'd21400: duty=88; 15'd21401: duty=101; 15'd21402: duty=114; 15'd21403: duty=104; 15'd21404: duty=110; 15'd21405: duty=104; 15'd21406: duty=103; 15'd21407: duty=111;
15'd21408: duty=108; 15'd21409: duty=110; 15'd21410: duty=103; 15'd21411: duty=100; 15'd21412: duty=101; 15'd21413: duty=108; 15'd21414: duty=96; 15'd21415: duty=90;
15'd21416: duty=84; 15'd21417: duty=90; 15'd21418: duty=98; 15'd21419: duty=101; 15'd21420: duty=108; 15'd21421: duty=106; 15'd21422: duty=121; 15'd21423: duty=116;
15'd21424: duty=121; 15'd21425: duty=125; 15'd21426: duty=125; 15'd21427: duty=124; 15'd21428: duty=137; 15'd21429: duty=133; 15'd21430: duty=127; 15'd21431: duty=139;
15'd21432: duty=131; 15'd21433: duty=129; 15'd21434: duty=131; 15'd21435: duty=145; 15'd21436: duty=157; 15'd21437: duty=163; 15'd21438: duty=165; 15'd21439: duty=176;
15'd21440: duty=168; 15'd21441: duty=164; 15'd21442: duty=163; 15'd21443: duty=165; 15'd21444: duty=168; 15'd21445: duty=167; 15'd21446: duty=171; 15'd21447: duty=160;
15'd21448: duty=166; 15'd21449: duty=161; 15'd21450: duty=167; 15'd21451: duty=159; 15'd21452: duty=166; 15'd21453: duty=167; 15'd21454: duty=172; 15'd21455: duty=171;
15'd21456: duty=165; 15'd21457: duty=166; 15'd21458: duty=149; 15'd21459: duty=146; 15'd21460: duty=145; 15'd21461: duty=142; 15'd21462: duty=138; 15'd21463: duty=134;
15'd21464: duty=131; 15'd21465: duty=139; 15'd21466: duty=140; 15'd21467: duty=136; 15'd21468: duty=132; 15'd21469: duty=133; 15'd21470: duty=127; 15'd21471: duty=122;
15'd21472: duty=121; 15'd21473: duty=128; 15'd21474: duty=123; 15'd21475: duty=115; 15'd21476: duty=107; 15'd21477: duty=92; 15'd21478: duty=92; 15'd21479: duty=109;
15'd21480: duty=104; 15'd21481: duty=95; 15'd21482: duty=96; 15'd21483: duty=99; 15'd21484: duty=105; 15'd21485: duty=91; 15'd21486: duty=102; 15'd21487: duty=109;
15'd21488: duty=96; 15'd21489: duty=100; 15'd21490: duty=95; 15'd21491: duty=94; 15'd21492: duty=93; 15'd21493: duty=87; 15'd21494: duty=102; 15'd21495: duty=106;
15'd21496: duty=96; 15'd21497: duty=109; 15'd21498: duty=118; 15'd21499: duty=115; 15'd21500: duty=111; 15'd21501: duty=112; 15'd21502: duty=106; 15'd21503: duty=116;
15'd21504: duty=113; 15'd21505: duty=118; 15'd21506: duty=128; 15'd21507: duty=126; 15'd21508: duty=142; 15'd21509: duty=130; 15'd21510: duty=136; 15'd21511: duty=131;
15'd21512: duty=135; 15'd21513: duty=139; 15'd21514: duty=142; 15'd21515: duty=135; 15'd21516: duty=155; 15'd21517: duty=169; 15'd21518: duty=163; 15'd21519: duty=176;
15'd21520: duty=169; 15'd21521: duty=160; 15'd21522: duty=163; 15'd21523: duty=168; 15'd21524: duty=161; 15'd21525: duty=164; 15'd21526: duty=166; 15'd21527: duty=167;
15'd21528: duty=157; 15'd21529: duty=148; 15'd21530: duty=153; 15'd21531: duty=164; 15'd21532: duty=165; 15'd21533: duty=165; 15'd21534: duty=153; 15'd21535: duty=157;
15'd21536: duty=152; 15'd21537: duty=145; 15'd21538: duty=142; 15'd21539: duty=139; 15'd21540: duty=144; 15'd21541: duty=135; 15'd21542: duty=137; 15'd21543: duty=140;
15'd21544: duty=134; 15'd21545: duty=130; 15'd21546: duty=132; 15'd21547: duty=128; 15'd21548: duty=123; 15'd21549: duty=126; 15'd21550: duty=125; 15'd21551: duty=111;
15'd21552: duty=112; 15'd21553: duty=114; 15'd21554: duty=100; 15'd21555: duty=115; 15'd21556: duty=113; 15'd21557: duty=105; 15'd21558: duty=118; 15'd21559: duty=114;
15'd21560: duty=106; 15'd21561: duty=105; 15'd21562: duty=97; 15'd21563: duty=107; 15'd21564: duty=100; 15'd21565: duty=94; 15'd21566: duty=110; 15'd21567: duty=109;
15'd21568: duty=114; 15'd21569: duty=104; 15'd21570: duty=95; 15'd21571: duty=99; 15'd21572: duty=102; 15'd21573: duty=102; 15'd21574: duty=115; 15'd21575: duty=118;
15'd21576: duty=123; 15'd21577: duty=127; 15'd21578: duty=119; 15'd21579: duty=110; 15'd21580: duty=115; 15'd21581: duty=128; 15'd21582: duty=131; 15'd21583: duty=122;
15'd21584: duty=123; 15'd21585: duty=129; 15'd21586: duty=135; 15'd21587: duty=135; 15'd21588: duty=136; 15'd21589: duty=137; 15'd21590: duty=135; 15'd21591: duty=142;
15'd21592: duty=142; 15'd21593: duty=140; 15'd21594: duty=153; 15'd21595: duty=157; 15'd21596: duty=157; 15'd21597: duty=159; 15'd21598: duty=159; 15'd21599: duty=177;
15'd21600: duty=170; 15'd21601: duty=163; 15'd21602: duty=164; 15'd21603: duty=157; 15'd21604: duty=159; 15'd21605: duty=161; 15'd21606: duty=154; 15'd21607: duty=154;
15'd21608: duty=148; 15'd21609: duty=160; 15'd21610: duty=159; 15'd21611: duty=153; 15'd21612: duty=150; 15'd21613: duty=150; 15'd21614: duty=147; 15'd21615: duty=151;
15'd21616: duty=145; 15'd21617: duty=140; 15'd21618: duty=133; 15'd21619: duty=127; 15'd21620: duty=134; 15'd21621: duty=131; 15'd21622: duty=132; 15'd21623: duty=125;
15'd21624: duty=125; 15'd21625: duty=125; 15'd21626: duty=132; 15'd21627: duty=116; 15'd21628: duty=121; 15'd21629: duty=118; 15'd21630: duty=108; 15'd21631: duty=113;
15'd21632: duty=118; 15'd21633: duty=118; 15'd21634: duty=110; 15'd21635: duty=101; 15'd21636: duty=103; 15'd21637: duty=114; 15'd21638: duty=111; 15'd21639: duty=110;
15'd21640: duty=105; 15'd21641: duty=96; 15'd21642: duty=108; 15'd21643: duty=109; 15'd21644: duty=106; 15'd21645: duty=98; 15'd21646: duty=101; 15'd21647: duty=101;
15'd21648: duty=94; 15'd21649: duty=102; 15'd21650: duty=107; 15'd21651: duty=112; 15'd21652: duty=105; 15'd21653: duty=107; 15'd21654: duty=106; 15'd21655: duty=110;
15'd21656: duty=113; 15'd21657: duty=113; 15'd21658: duty=130; 15'd21659: duty=126; 15'd21660: duty=115; 15'd21661: duty=119; 15'd21662: duty=127; 15'd21663: duty=131;
15'd21664: duty=128; 15'd21665: duty=131; 15'd21666: duty=133; 15'd21667: duty=137; 15'd21668: duty=136; 15'd21669: duty=142; 15'd21670: duty=150; 15'd21671: duty=151;
15'd21672: duty=147; 15'd21673: duty=158; 15'd21674: duty=165; 15'd21675: duty=168; 15'd21676: duty=179; 15'd21677: duty=170; 15'd21678: duty=173; 15'd21679: duty=174;
15'd21680: duty=168; 15'd21681: duty=171; 15'd21682: duty=160; 15'd21683: duty=163; 15'd21684: duty=160; 15'd21685: duty=159; 15'd21686: duty=155; 15'd21687: duty=145;
15'd21688: duty=140; 15'd21689: duty=146; 15'd21690: duty=150; 15'd21691: duty=149; 15'd21692: duty=160; 15'd21693: duty=159; 15'd21694: duty=158; 15'd21695: duty=147;
15'd21696: duty=153; 15'd21697: duty=144; 15'd21698: duty=142; 15'd21699: duty=140; 15'd21700: duty=129; 15'd21701: duty=117; 15'd21702: duty=117; 15'd21703: duty=114;
15'd21704: duty=120; 15'd21705: duty=126; 15'd21706: duty=115; 15'd21707: duty=116; 15'd21708: duty=106; 15'd21709: duty=117; 15'd21710: duty=115; 15'd21711: duty=119;
15'd21712: duty=112; 15'd21713: duty=100; 15'd21714: duty=112; 15'd21715: duty=98; 15'd21716: duty=98; 15'd21717: duty=99; 15'd21718: duty=93; 15'd21719: duty=93;
15'd21720: duty=100; 15'd21721: duty=108; 15'd21722: duty=109; 15'd21723: duty=107; 15'd21724: duty=100; 15'd21725: duty=104; 15'd21726: duty=102; 15'd21727: duty=104;
15'd21728: duty=110; 15'd21729: duty=104; 15'd21730: duty=121; 15'd21731: duty=121; 15'd21732: duty=104; 15'd21733: duty=109; 15'd21734: duty=115; 15'd21735: duty=122;
15'd21736: duty=120; 15'd21737: duty=131; 15'd21738: duty=133; 15'd21739: duty=134; 15'd21740: duty=132; 15'd21741: duty=125; 15'd21742: duty=130; 15'd21743: duty=120;
15'd21744: duty=126; 15'd21745: duty=134; 15'd21746: duty=135; 15'd21747: duty=138; 15'd21748: duty=140; 15'd21749: duty=150; 15'd21750: duty=158; 15'd21751: duty=162;
15'd21752: duty=169; 15'd21753: duty=168; 15'd21754: duty=158; 15'd21755: duty=159; 15'd21756: duty=172; 15'd21757: duty=157; 15'd21758: duty=155; 15'd21759: duty=153;
15'd21760: duty=137; 15'd21761: duty=146; 15'd21762: duty=157; 15'd21763: duty=160; 15'd21764: duty=160; 15'd21765: duty=156; 15'd21766: duty=153; 15'd21767: duty=151;
15'd21768: duty=160; 15'd21769: duty=158; 15'd21770: duty=156; 15'd21771: duty=162; 15'd21772: duty=152; 15'd21773: duty=145; 15'd21774: duty=146; 15'd21775: duty=144;
15'd21776: duty=142; 15'd21777: duty=136; 15'd21778: duty=137; 15'd21779: duty=152; 15'd21780: duty=152; 15'd21781: duty=138; 15'd21782: duty=128; 15'd21783: duty=109;
15'd21784: duty=114; 15'd21785: duty=118; 15'd21786: duty=100; 15'd21787: duty=95; 15'd21788: duty=89; 15'd21789: duty=101; 15'd21790: duty=112; 15'd21791: duty=105;
15'd21792: duty=94; 15'd21793: duty=98; 15'd21794: duty=105; 15'd21795: duty=100; 15'd21796: duty=110; 15'd21797: duty=111; 15'd21798: duty=109; 15'd21799: duty=91;
15'd21800: duty=98; 15'd21801: duty=104; 15'd21802: duty=96; 15'd21803: duty=100; 15'd21804: duty=91; 15'd21805: duty=108; 15'd21806: duty=97; 15'd21807: duty=102;
15'd21808: duty=117; 15'd21809: duty=116; 15'd21810: duty=128; 15'd21811: duty=135; 15'd21812: duty=132; 15'd21813: duty=125; 15'd21814: duty=127; 15'd21815: duty=123;
15'd21816: duty=114; 15'd21817: duty=117; 15'd21818: duty=137; 15'd21819: duty=141; 15'd21820: duty=139; 15'd21821: duty=144; 15'd21822: duty=143; 15'd21823: duty=133;
15'd21824: duty=140; 15'd21825: duty=145; 15'd21826: duty=143; 15'd21827: duty=145; 15'd21828: duty=151; 15'd21829: duty=165; 15'd21830: duty=162; 15'd21831: duty=158;
15'd21832: duty=157; 15'd21833: duty=159; 15'd21834: duty=159; 15'd21835: duty=157; 15'd21836: duty=159; 15'd21837: duty=159; 15'd21838: duty=164; 15'd21839: duty=167;
15'd21840: duty=160; 15'd21841: duty=151; 15'd21842: duty=148; 15'd21843: duty=151; 15'd21844: duty=151; 15'd21845: duty=150; 15'd21846: duty=153; 15'd21847: duty=154;
15'd21848: duty=148; 15'd21849: duty=139; 15'd21850: duty=136; 15'd21851: duty=140; 15'd21852: duty=137; 15'd21853: duty=139; 15'd21854: duty=139; 15'd21855: duty=131;
15'd21856: duty=119; 15'd21857: duty=119; 15'd21858: duty=118; 15'd21859: duty=134; 15'd21860: duty=136; 15'd21861: duty=130; 15'd21862: duty=126; 15'd21863: duty=118;
15'd21864: duty=126; 15'd21865: duty=117; 15'd21866: duty=112; 15'd21867: duty=105; 15'd21868: duty=104; 15'd21869: duty=99; 15'd21870: duty=110; 15'd21871: duty=108;
15'd21872: duty=101; 15'd21873: duty=99; 15'd21874: duty=102; 15'd21875: duty=110; 15'd21876: duty=110; 15'd21877: duty=107; 15'd21878: duty=105; 15'd21879: duty=104;
15'd21880: duty=99; 15'd21881: duty=106; 15'd21882: duty=98; 15'd21883: duty=100; 15'd21884: duty=107; 15'd21885: duty=104; 15'd21886: duty=116; 15'd21887: duty=123;
15'd21888: duty=111; 15'd21889: duty=115; 15'd21890: duty=108; 15'd21891: duty=113; 15'd21892: duty=127; 15'd21893: duty=126; 15'd21894: duty=124; 15'd21895: duty=130;
15'd21896: duty=128; 15'd21897: duty=139; 15'd21898: duty=143; 15'd21899: duty=139; 15'd21900: duty=149; 15'd21901: duty=141; 15'd21902: duty=144; 15'd21903: duty=144;
15'd21904: duty=141; 15'd21905: duty=149; 15'd21906: duty=159; 15'd21907: duty=158; 15'd21908: duty=161; 15'd21909: duty=169; 15'd21910: duty=172; 15'd21911: duty=176;
15'd21912: duty=166; 15'd21913: duty=158; 15'd21914: duty=152; 15'd21915: duty=151; 15'd21916: duty=149; 15'd21917: duty=146; 15'd21918: duty=149; 15'd21919: duty=142;
15'd21920: duty=154; 15'd21921: duty=153; 15'd21922: duty=160; 15'd21923: duty=161; 15'd21924: duty=149; 15'd21925: duty=148; 15'd21926: duty=151; 15'd21927: duty=154;
15'd21928: duty=145; 15'd21929: duty=138; 15'd21930: duty=132; 15'd21931: duty=133; 15'd21932: duty=132; 15'd21933: duty=125; 15'd21934: duty=127; 15'd21935: duty=127;
15'd21936: duty=122; 15'd21937: duty=125; 15'd21938: duty=122; 15'd21939: duty=122; 15'd21940: duty=124; 15'd21941: duty=122; 15'd21942: duty=109; 15'd21943: duty=107;
15'd21944: duty=113; 15'd21945: duty=104; 15'd21946: duty=106; 15'd21947: duty=110; 15'd21948: duty=102; 15'd21949: duty=110; 15'd21950: duty=104; 15'd21951: duty=110;
15'd21952: duty=104; 15'd21953: duty=104; 15'd21954: duty=115; 15'd21955: duty=99; 15'd21956: duty=110; 15'd21957: duty=111; 15'd21958: duty=107; 15'd21959: duty=102;
15'd21960: duty=103; 15'd21961: duty=108; 15'd21962: duty=110; 15'd21963: duty=118; 15'd21964: duty=112; 15'd21965: duty=119; 15'd21966: duty=121; 15'd21967: duty=125;
15'd21968: duty=122; 15'd21969: duty=123; 15'd21970: duty=126; 15'd21971: duty=125; 15'd21972: duty=133; 15'd21973: duty=125; 15'd21974: duty=130; 15'd21975: duty=132;
15'd21976: duty=135; 15'd21977: duty=145; 15'd21978: duty=139; 15'd21979: duty=140; 15'd21980: duty=138; 15'd21981: duty=137; 15'd21982: duty=146; 15'd21983: duty=138;
15'd21984: duty=148; 15'd21985: duty=163; 15'd21986: duty=173; 15'd21987: duty=169; 15'd21988: duty=167; 15'd21989: duty=166; 15'd21990: duty=167; 15'd21991: duty=172;
15'd21992: duty=160; 15'd21993: duty=166; 15'd21994: duty=166; 15'd21995: duty=168; 15'd21996: duty=165; 15'd21997: duty=151; 15'd21998: duty=148; 15'd21999: duty=150;
15'd22000: duty=155; 15'd22001: duty=159; 15'd22002: duty=157; 15'd22003: duty=158; 15'd22004: duty=157; 15'd22005: duty=148; 15'd22006: duty=151; 15'd22007: duty=146;
15'd22008: duty=127; 15'd22009: duty=127; 15'd22010: duty=121; 15'd22011: duty=122; 15'd22012: duty=124; 15'd22013: duty=124; 15'd22014: duty=123; 15'd22015: duty=117;
15'd22016: duty=115; 15'd22017: duty=112; 15'd22018: duty=116; 15'd22019: duty=112; 15'd22020: duty=120; 15'd22021: duty=113; 15'd22022: duty=110; 15'd22023: duty=105;
15'd22024: duty=93; 15'd22025: duty=95; 15'd22026: duty=90; 15'd22027: duty=99; 15'd22028: duty=93; 15'd22029: duty=104; 15'd22030: duty=111; 15'd22031: duty=107;
15'd22032: duty=114; 15'd22033: duty=107; 15'd22034: duty=108; 15'd22035: duty=99; 15'd22036: duty=90; 15'd22037: duty=96; 15'd22038: duty=109; 15'd22039: duty=110;
15'd22040: duty=107; 15'd22041: duty=102; 15'd22042: duty=106; 15'd22043: duty=111; 15'd22044: duty=104; 15'd22045: duty=118; 15'd22046: duty=123; 15'd22047: duty=125;
15'd22048: duty=131; 15'd22049: duty=119; 15'd22050: duty=123; 15'd22051: duty=124; 15'd22052: duty=119; 15'd22053: duty=128; 15'd22054: duty=124; 15'd22055: duty=125;
15'd22056: duty=136; 15'd22057: duty=137; 15'd22058: duty=131; 15'd22059: duty=142; 15'd22060: duty=152; 15'd22061: duty=145; 15'd22062: duty=156; 15'd22063: duty=157;
15'd22064: duty=157; 15'd22065: duty=168; 15'd22066: duty=174; 15'd22067: duty=176; 15'd22068: duty=171; 15'd22069: duty=165; 15'd22070: duty=158; 15'd22071: duty=159;
15'd22072: duty=153; 15'd22073: duty=157; 15'd22074: duty=163; 15'd22075: duty=164; 15'd22076: duty=163; 15'd22077: duty=163; 15'd22078: duty=169; 15'd22079: duty=173;
15'd22080: duty=179; 15'd22081: duty=173; 15'd22082: duty=174; 15'd22083: duty=161; 15'd22084: duty=148; 15'd22085: duty=145; 15'd22086: duty=143; 15'd22087: duty=157;
15'd22088: duty=149; 15'd22089: duty=136; 15'd22090: duty=134; 15'd22091: duty=137; 15'd22092: duty=135; 15'd22093: duty=126; 15'd22094: duty=142; 15'd22095: duty=126;
15'd22096: duty=108; 15'd22097: duty=112; 15'd22098: duty=114; 15'd22099: duty=118; 15'd22100: duty=109; 15'd22101: duty=98; 15'd22102: duty=69; 15'd22103: duty=81;
15'd22104: duty=99; 15'd22105: duty=110; 15'd22106: duty=105; 15'd22107: duty=107; 15'd22108: duty=99; 15'd22109: duty=87; 15'd22110: duty=88; 15'd22111: duty=80;
15'd22112: duty=87; 15'd22113: duty=85; 15'd22114: duty=85; 15'd22115: duty=87; 15'd22116: duty=97; 15'd22117: duty=104; 15'd22118: duty=104; 15'd22119: duty=101;
15'd22120: duty=111; 15'd22121: duty=112; 15'd22122: duty=120; 15'd22123: duty=115; 15'd22124: duty=119; 15'd22125: duty=121; 15'd22126: duty=117; 15'd22127: duty=118;
15'd22128: duty=129; 15'd22129: duty=129; 15'd22130: duty=121; 15'd22131: duty=134; 15'd22132: duty=131; 15'd22133: duty=129; 15'd22134: duty=139; 15'd22135: duty=133;
15'd22136: duty=148; 15'd22137: duty=149; 15'd22138: duty=139; 15'd22139: duty=152; 15'd22140: duty=149; 15'd22141: duty=155; 15'd22142: duty=159; 15'd22143: duty=159;
15'd22144: duty=160; 15'd22145: duty=172; 15'd22146: duty=163; 15'd22147: duty=172; 15'd22148: duty=171; 15'd22149: duty=161; 15'd22150: duty=163; 15'd22151: duty=158;
15'd22152: duty=157; 15'd22153: duty=165; 15'd22154: duty=157; 15'd22155: duty=155; 15'd22156: duty=154; 15'd22157: duty=162; 15'd22158: duty=166; 15'd22159: duty=157;
15'd22160: duty=163; 15'd22161: duty=163; 15'd22162: duty=163; 15'd22163: duty=155; 15'd22164: duty=155; 15'd22165: duty=142; 15'd22166: duty=134; 15'd22167: duty=135;
15'd22168: duty=140; 15'd22169: duty=135; 15'd22170: duty=137; 15'd22171: duty=133; 15'd22172: duty=124; 15'd22173: duty=118; 15'd22174: duty=116; 15'd22175: duty=114;
15'd22176: duty=122; 15'd22177: duty=118; 15'd22178: duty=109; 15'd22179: duty=106; 15'd22180: duty=96; 15'd22181: duty=96; 15'd22182: duty=102; 15'd22183: duty=98;
15'd22184: duty=103; 15'd22185: duty=103; 15'd22186: duty=94; 15'd22187: duty=95; 15'd22188: duty=80; 15'd22189: duty=86; 15'd22190: duty=90; 15'd22191: duty=95;
15'd22192: duty=82; 15'd22193: duty=79; 15'd22194: duty=90; 15'd22195: duty=100; 15'd22196: duty=122; 15'd22197: duty=109; 15'd22198: duty=110; 15'd22199: duty=112;
15'd22200: duty=109; 15'd22201: duty=116; 15'd22202: duty=110; 15'd22203: duty=101; 15'd22204: duty=102; 15'd22205: duty=108; 15'd22206: duty=121; 15'd22207: duty=131;
15'd22208: duty=124; 15'd22209: duty=124; 15'd22210: duty=128; 15'd22211: duty=137; 15'd22212: duty=140; 15'd22213: duty=137; 15'd22214: duty=138; 15'd22215: duty=148;
15'd22216: duty=153; 15'd22217: duty=145; 15'd22218: duty=147; 15'd22219: duty=160; 15'd22220: duty=167; 15'd22221: duty=169; 15'd22222: duty=173; 15'd22223: duty=189;
15'd22224: duty=181; 15'd22225: duty=182; 15'd22226: duty=183; 15'd22227: duty=182; 15'd22228: duty=178; 15'd22229: duty=166; 15'd22230: duty=167; 15'd22231: duty=161;
15'd22232: duty=159; 15'd22233: duty=152; 15'd22234: duty=158; 15'd22235: duty=160; 15'd22236: duty=153; 15'd22237: duty=151; 15'd22238: duty=157; 15'd22239: duty=165;
15'd22240: duty=153; 15'd22241: duty=151; 15'd22242: duty=154; 15'd22243: duty=141; 15'd22244: duty=137; 15'd22245: duty=136; 15'd22246: duty=130; 15'd22247: duty=134;
15'd22248: duty=128; 15'd22249: duty=119; 15'd22250: duty=122; 15'd22251: duty=110; 15'd22252: duty=119; 15'd22253: duty=114; 15'd22254: duty=114; 15'd22255: duty=115;
15'd22256: duty=102; 15'd22257: duty=98; 15'd22258: duty=94; 15'd22259: duty=106; 15'd22260: duty=107; 15'd22261: duty=104; 15'd22262: duty=97; 15'd22263: duty=111;
15'd22264: duty=105; 15'd22265: duty=104; 15'd22266: duty=104; 15'd22267: duty=106; 15'd22268: duty=97; 15'd22269: duty=78; 15'd22270: duty=77; 15'd22271: duty=80;
15'd22272: duty=92; 15'd22273: duty=94; 15'd22274: duty=104; 15'd22275: duty=93; 15'd22276: duty=99; 15'd22277: duty=112; 15'd22278: duty=113; 15'd22279: duty=119;
15'd22280: duty=117; 15'd22281: duty=119; 15'd22282: duty=128; 15'd22283: duty=130; 15'd22284: duty=122; 15'd22285: duty=130; 15'd22286: duty=122; 15'd22287: duty=119;
15'd22288: duty=106; 15'd22289: duty=112; 15'd22290: duty=135; 15'd22291: duty=137; 15'd22292: duty=134; 15'd22293: duty=134; 15'd22294: duty=133; 15'd22295: duty=144;
15'd22296: duty=168; 15'd22297: duty=166; 15'd22298: duty=161; 15'd22299: duty=172; 15'd22300: duty=168; 15'd22301: duty=170; 15'd22302: duty=187; 15'd22303: duty=172;
15'd22304: duty=173; 15'd22305: duty=162; 15'd22306: duty=152; 15'd22307: duty=158; 15'd22308: duty=152; 15'd22309: duty=152; 15'd22310: duty=164; 15'd22311: duty=163;
15'd22312: duty=157; 15'd22313: duty=169; 15'd22314: duty=169; 15'd22315: duty=167; 15'd22316: duty=165; 15'd22317: duty=156; 15'd22318: duty=162; 15'd22319: duty=165;
15'd22320: duty=159; 15'd22321: duty=153; 15'd22322: duty=152; 15'd22323: duty=140; 15'd22324: duty=136; 15'd22325: duty=120; 15'd22326: duty=121; 15'd22327: duty=123;
15'd22328: duty=124; 15'd22329: duty=127; 15'd22330: duty=121; 15'd22331: duty=122; 15'd22332: duty=119; 15'd22333: duty=119; 15'd22334: duty=106; 15'd22335: duty=118;
15'd22336: duty=115; 15'd22337: duty=105; 15'd22338: duty=103; 15'd22339: duty=97; 15'd22340: duty=98; 15'd22341: duty=105; 15'd22342: duty=99; 15'd22343: duty=101;
15'd22344: duty=98; 15'd22345: duty=101; 15'd22346: duty=90; 15'd22347: duty=96; 15'd22348: duty=104; 15'd22349: duty=104; 15'd22350: duty=110; 15'd22351: duty=91;
15'd22352: duty=95; 15'd22353: duty=104; 15'd22354: duty=110; 15'd22355: duty=104; 15'd22356: duty=110; 15'd22357: duty=122; 15'd22358: duty=115; 15'd22359: duty=122;
15'd22360: duty=105; 15'd22361: duty=102; 15'd22362: duty=118; 15'd22363: duty=114; 15'd22364: duty=127; 15'd22365: duty=121; 15'd22366: duty=126; 15'd22367: duty=122;
15'd22368: duty=126; 15'd22369: duty=117; 15'd22370: duty=136; 15'd22371: duty=131; 15'd22372: duty=124; 15'd22373: duty=137; 15'd22374: duty=130; 15'd22375: duty=161;
15'd22376: duty=170; 15'd22377: duty=170; 15'd22378: duty=161; 15'd22379: duty=169; 15'd22380: duty=161; 15'd22381: duty=154; 15'd22382: duty=164; 15'd22383: duty=151;
15'd22384: duty=148; 15'd22385: duty=155; 15'd22386: duty=161; 15'd22387: duty=162; 15'd22388: duty=176; 15'd22389: duty=177; 15'd22390: duty=177; 15'd22391: duty=170;
15'd22392: duty=173; 15'd22393: duty=167; 15'd22394: duty=164; 15'd22395: duty=172; 15'd22396: duty=161; 15'd22397: duty=155; 15'd22398: duty=146; 15'd22399: duty=147;
15'd22400: duty=136; 15'd22401: duty=141; 15'd22402: duty=141; 15'd22403: duty=129; 15'd22404: duty=131; 15'd22405: duty=139; 15'd22406: duty=128; 15'd22407: duty=126;
15'd22408: duty=129; 15'd22409: duty=120; 15'd22410: duty=113; 15'd22411: duty=112; 15'd22412: duty=102; 15'd22413: duty=103; 15'd22414: duty=100; 15'd22415: duty=103;
15'd22416: duty=110; 15'd22417: duty=99; 15'd22418: duty=106; 15'd22419: duty=103; 15'd22420: duty=86; 15'd22421: duty=91; 15'd22422: duty=108; 15'd22423: duty=102;
15'd22424: duty=101; 15'd22425: duty=94; 15'd22426: duty=98; 15'd22427: duty=94; 15'd22428: duty=80; 15'd22429: duty=102; 15'd22430: duty=123; 15'd22431: duty=113;
15'd22432: duty=114; 15'd22433: duty=102; 15'd22434: duty=106; 15'd22435: duty=110; 15'd22436: duty=110; 15'd22437: duty=116; 15'd22438: duty=121; 15'd22439: duty=115;
15'd22440: duty=113; 15'd22441: duty=124; 15'd22442: duty=124; 15'd22443: duty=127; 15'd22444: duty=128; 15'd22445: duty=137; 15'd22446: duty=146; 15'd22447: duty=138;
15'd22448: duty=140; 15'd22449: duty=140; 15'd22450: duty=131; 15'd22451: duty=131; 15'd22452: duty=136; 15'd22453: duty=158; 15'd22454: duty=171; 15'd22455: duty=162;
15'd22456: duty=157; 15'd22457: duty=164; 15'd22458: duty=168; 15'd22459: duty=163; 15'd22460: duty=154; 15'd22461: duty=160; 15'd22462: duty=168; 15'd22463: duty=159;
15'd22464: duty=150; 15'd22465: duty=145; 15'd22466: duty=134; 15'd22467: duty=145; 15'd22468: duty=153; 15'd22469: duty=162; 15'd22470: duty=159; 15'd22471: duty=163;
15'd22472: duty=162; 15'd22473: duty=157; 15'd22474: duty=147; 15'd22475: duty=149; 15'd22476: duty=150; 15'd22477: duty=138; 15'd22478: duty=136; 15'd22479: duty=128;
15'd22480: duty=135; 15'd22481: duty=135; 15'd22482: duty=126; 15'd22483: duty=123; 15'd22484: duty=129; 15'd22485: duty=126; 15'd22486: duty=122; 15'd22487: duty=125;
15'd22488: duty=127; 15'd22489: duty=120; 15'd22490: duty=109; 15'd22491: duty=112; 15'd22492: duty=115; 15'd22493: duty=102; 15'd22494: duty=107; 15'd22495: duty=114;
15'd22496: duty=105; 15'd22497: duty=96; 15'd22498: duty=100; 15'd22499: duty=111; 15'd22500: duty=106; 15'd22501: duty=106; 15'd22502: duty=112; 15'd22503: duty=116;
15'd22504: duty=118; 15'd22505: duty=106; 15'd22506: duty=106; 15'd22507: duty=97; 15'd22508: duty=101; 15'd22509: duty=103; 15'd22510: duty=107; 15'd22511: duty=117;
15'd22512: duty=111; 15'd22513: duty=117; 15'd22514: duty=118; 15'd22515: duty=123; 15'd22516: duty=124; 15'd22517: duty=129; 15'd22518: duty=134; 15'd22519: duty=138;
15'd22520: duty=141; 15'd22521: duty=137; 15'd22522: duty=133; 15'd22523: duty=137; 15'd22524: duty=132; 15'd22525: duty=128; 15'd22526: duty=118; 15'd22527: duty=131;
15'd22528: duty=135; 15'd22529: duty=142; 15'd22530: duty=158; 15'd22531: duty=171; 15'd22532: duty=181; 15'd22533: duty=163; 15'd22534: duty=164; 15'd22535: duty=152;
15'd22536: duty=150; 15'd22537: duty=157; 15'd22538: duty=158; 15'd22539: duty=157; 15'd22540: duty=142; 15'd22541: duty=139; 15'd22542: duty=137; 15'd22543: duty=142;
15'd22544: duty=155; 15'd22545: duty=148; 15'd22546: duty=150; 15'd22547: duty=154; 15'd22548: duty=159; 15'd22549: duty=159; 15'd22550: duty=160; 15'd22551: duty=152;
15'd22552: duty=145; 15'd22553: duty=134; 15'd22554: duty=134; 15'd22555: duty=140; 15'd22556: duty=134; 15'd22557: duty=128; 15'd22558: duty=125; 15'd22559: duty=134;
15'd22560: duty=128; 15'd22561: duty=142; 15'd22562: duty=140; 15'd22563: duty=130; 15'd22564: duty=110; 15'd22565: duty=99; 15'd22566: duty=105; 15'd22567: duty=112;
15'd22568: duty=114; 15'd22569: duty=109; 15'd22570: duty=102; 15'd22571: duty=96; 15'd22572: duty=102; 15'd22573: duty=98; 15'd22574: duty=118; 15'd22575: duty=115;
15'd22576: duty=105; 15'd22577: duty=107; 15'd22578: duty=116; 15'd22579: duty=115; 15'd22580: duty=108; 15'd22581: duty=93; 15'd22582: duty=81; 15'd22583: duty=87;
15'd22584: duty=97; 15'd22585: duty=118; 15'd22586: duty=116; 15'd22587: duty=112; 15'd22588: duty=108; 15'd22589: duty=110; 15'd22590: duty=120; 15'd22591: duty=127;
15'd22592: duty=127; 15'd22593: duty=115; 15'd22594: duty=122; 15'd22595: duty=126; 15'd22596: duty=124; 15'd22597: duty=124; 15'd22598: duty=127; 15'd22599: duty=120;
15'd22600: duty=122; 15'd22601: duty=127; 15'd22602: duty=131; 15'd22603: duty=142; 15'd22604: duty=153; 15'd22605: duty=158; 15'd22606: duty=151; 15'd22607: duty=153;
15'd22608: duty=150; 15'd22609: duty=145; 15'd22610: duty=149; 15'd22611: duty=160; 15'd22612: duty=165; 15'd22613: duty=164; 15'd22614: duty=167; 15'd22615: duty=170;
15'd22616: duty=167; 15'd22617: duty=162; 15'd22618: duty=161; 15'd22619: duty=165; 15'd22620: duty=160; 15'd22621: duty=154; 15'd22622: duty=160; 15'd22623: duty=163;
15'd22624: duty=150; 15'd22625: duty=153; 15'd22626: duty=162; 15'd22627: duty=157; 15'd22628: duty=148; 15'd22629: duty=148; 15'd22630: duty=147; 15'd22631: duty=132;
15'd22632: duty=134; 15'd22633: duty=140; 15'd22634: duty=148; 15'd22635: duty=139; 15'd22636: duty=127; 15'd22637: duty=130; 15'd22638: duty=124; 15'd22639: duty=116;
15'd22640: duty=116; 15'd22641: duty=116; 15'd22642: duty=119; 15'd22643: duty=116; 15'd22644: duty=123; 15'd22645: duty=121; 15'd22646: duty=110; 15'd22647: duty=114;
15'd22648: duty=112; 15'd22649: duty=106; 15'd22650: duty=96; 15'd22651: duty=95; 15'd22652: duty=98; 15'd22653: duty=99; 15'd22654: duty=104; 15'd22655: duty=100;
15'd22656: duty=107; 15'd22657: duty=111; 15'd22658: duty=100; 15'd22659: duty=100; 15'd22660: duty=106; 15'd22661: duty=118; 15'd22662: duty=114; 15'd22663: duty=116;
15'd22664: duty=119; 15'd22665: duty=113; 15'd22666: duty=112; 15'd22667: duty=115; 15'd22668: duty=112; 15'd22669: duty=109; 15'd22670: duty=118; 15'd22671: duty=113;
15'd22672: duty=117; 15'd22673: duty=119; 15'd22674: duty=123; 15'd22675: duty=137; 15'd22676: duty=129; 15'd22677: duty=131; 15'd22678: duty=136; 15'd22679: duty=128;
15'd22680: duty=126; 15'd22681: duty=134; 15'd22682: duty=133; 15'd22683: duty=132; 15'd22684: duty=138; 15'd22685: duty=142; 15'd22686: duty=159; 15'd22687: duty=163;
15'd22688: duty=157; 15'd22689: duty=160; 15'd22690: duty=156; 15'd22691: duty=150; 15'd22692: duty=155; 15'd22693: duty=149; 15'd22694: duty=149; 15'd22695: duty=149;
15'd22696: duty=154; 15'd22697: duty=157; 15'd22698: duty=160; 15'd22699: duty=156; 15'd22700: duty=157; 15'd22701: duty=162; 15'd22702: duty=152; 15'd22703: duty=151;
15'd22704: duty=157; 15'd22705: duty=153; 15'd22706: duty=140; 15'd22707: duty=147; 15'd22708: duty=149; 15'd22709: duty=142; 15'd22710: duty=137; 15'd22711: duty=145;
15'd22712: duty=142; 15'd22713: duty=133; 15'd22714: duty=137; 15'd22715: duty=131; 15'd22716: duty=131; 15'd22717: duty=129; 15'd22718: duty=128; 15'd22719: duty=130;
15'd22720: duty=118; 15'd22721: duty=104; 15'd22722: duty=107; 15'd22723: duty=110; 15'd22724: duty=109; 15'd22725: duty=105; 15'd22726: duty=112; 15'd22727: duty=104;
15'd22728: duty=93; 15'd22729: duty=94; 15'd22730: duty=95; 15'd22731: duty=105; 15'd22732: duty=104; 15'd22733: duty=114; 15'd22734: duty=118; 15'd22735: duty=118;
15'd22736: duty=112; 15'd22737: duty=117; 15'd22738: duty=111; 15'd22739: duty=96; 15'd22740: duty=95; 15'd22741: duty=101; 15'd22742: duty=123; 15'd22743: duty=121;
15'd22744: duty=127; 15'd22745: duty=121; 15'd22746: duty=121; 15'd22747: duty=127; 15'd22748: duty=126; 15'd22749: duty=134; 15'd22750: duty=142; 15'd22751: duty=145;
15'd22752: duty=148; 15'd22753: duty=134; 15'd22754: duty=130; 15'd22755: duty=146; 15'd22756: duty=139; 15'd22757: duty=130; 15'd22758: duty=132; 15'd22759: duty=135;
15'd22760: duty=143; 15'd22761: duty=151; 15'd22762: duty=142; 15'd22763: duty=151; 15'd22764: duty=145; 15'd22765: duty=138; 15'd22766: duty=148; 15'd22767: duty=154;
15'd22768: duty=168; 15'd22769: duty=166; 15'd22770: duty=161; 15'd22771: duty=158; 15'd22772: duty=154; 15'd22773: duty=149; 15'd22774: duty=156; 15'd22775: duty=144;
15'd22776: duty=137; 15'd22777: duty=142; 15'd22778: duty=155; 15'd22779: duty=163; 15'd22780: duty=162; 15'd22781: duty=157; 15'd22782: duty=145; 15'd22783: duty=135;
15'd22784: duty=135; 15'd22785: duty=135; 15'd22786: duty=125; 15'd22787: duty=129; 15'd22788: duty=133; 15'd22789: duty=132; 15'd22790: duty=122; 15'd22791: duty=130;
15'd22792: duty=123; 15'd22793: duty=121; 15'd22794: duty=116; 15'd22795: duty=125; 15'd22796: duty=132; 15'd22797: duty=124; 15'd22798: duty=122; 15'd22799: duty=107;
15'd22800: duty=107; 15'd22801: duty=101; 15'd22802: duty=99; 15'd22803: duty=112; 15'd22804: duty=106; 15'd22805: duty=103; 15'd22806: duty=106; 15'd22807: duty=109;
15'd22808: duty=123; 15'd22809: duty=115; 15'd22810: duty=117; 15'd22811: duty=115; 15'd22812: duty=110; 15'd22813: duty=109; 15'd22814: duty=102; 15'd22815: duty=97;
15'd22816: duty=93; 15'd22817: duty=100; 15'd22818: duty=106; 15'd22819: duty=109; 15'd22820: duty=105; 15'd22821: duty=109; 15'd22822: duty=117; 15'd22823: duty=115;
15'd22824: duty=134; 15'd22825: duty=130; 15'd22826: duty=135; 15'd22827: duty=133; 15'd22828: duty=129; 15'd22829: duty=128; 15'd22830: duty=129; 15'd22831: duty=131;
15'd22832: duty=126; 15'd22833: duty=130; 15'd22834: duty=133; 15'd22835: duty=141; 15'd22836: duty=138; 15'd22837: duty=149; 15'd22838: duty=149; 15'd22839: duty=160;
15'd22840: duty=158; 15'd22841: duty=158; 15'd22842: duty=170; 15'd22843: duty=165; 15'd22844: duty=168; 15'd22845: duty=169; 15'd22846: duty=162; 15'd22847: duty=160;
15'd22848: duty=154; 15'd22849: duty=145; 15'd22850: duty=151; 15'd22851: duty=156; 15'd22852: duty=154; 15'd22853: duty=165; 15'd22854: duty=161; 15'd22855: duty=157;
15'd22856: duty=157; 15'd22857: duty=149; 15'd22858: duty=152; 15'd22859: duty=152; 15'd22860: duty=145; 15'd22861: duty=137; 15'd22862: duty=140; 15'd22863: duty=136;
15'd22864: duty=131; 15'd22865: duty=133; 15'd22866: duty=130; 15'd22867: duty=136; 15'd22868: duty=131; 15'd22869: duty=128; 15'd22870: duty=128; 15'd22871: duty=125;
15'd22872: duty=124; 15'd22873: duty=118; 15'd22874: duty=116; 15'd22875: duty=109; 15'd22876: duty=110; 15'd22877: duty=108; 15'd22878: duty=112; 15'd22879: duty=108;
15'd22880: duty=101; 15'd22881: duty=102; 15'd22882: duty=101; 15'd22883: duty=108; 15'd22884: duty=110; 15'd22885: duty=107; 15'd22886: duty=95; 15'd22887: duty=101;
15'd22888: duty=104; 15'd22889: duty=103; 15'd22890: duty=115; 15'd22891: duty=94; 15'd22892: duty=90; 15'd22893: duty=84; 15'd22894: duty=98; 15'd22895: duty=113;
15'd22896: duty=115; 15'd22897: duty=121; 15'd22898: duty=115; 15'd22899: duty=126; 15'd22900: duty=134; 15'd22901: duty=129; 15'd22902: duty=121; 15'd22903: duty=129;
15'd22904: duty=124; 15'd22905: duty=134; 15'd22906: duty=139; 15'd22907: duty=136; 15'd22908: duty=133; 15'd22909: duty=131; 15'd22910: duty=139; 15'd22911: duty=148;
15'd22912: duty=144; 15'd22913: duty=142; 15'd22914: duty=144; 15'd22915: duty=140; 15'd22916: duty=150; 15'd22917: duty=153; 15'd22918: duty=153; 15'd22919: duty=157;
15'd22920: duty=153; 15'd22921: duty=157; 15'd22922: duty=158; 15'd22923: duty=164; 15'd22924: duty=170; 15'd22925: duty=158; 15'd22926: duty=157; 15'd22927: duty=154;
15'd22928: duty=152; 15'd22929: duty=155; 15'd22930: duty=154; 15'd22931: duty=154; 15'd22932: duty=148; 15'd22933: duty=152; 15'd22934: duty=152; 15'd22935: duty=149;
15'd22936: duty=151; 15'd22937: duty=152; 15'd22938: duty=153; 15'd22939: duty=148; 15'd22940: duty=148; 15'd22941: duty=145; 15'd22942: duty=137; 15'd22943: duty=127;
15'd22944: duty=124; 15'd22945: duty=129; 15'd22946: duty=120; 15'd22947: duty=118; 15'd22948: duty=123; 15'd22949: duty=120; 15'd22950: duty=121; 15'd22951: duty=113;
15'd22952: duty=120; 15'd22953: duty=112; 15'd22954: duty=107; 15'd22955: duty=106; 15'd22956: duty=99; 15'd22957: duty=110; 15'd22958: duty=96; 15'd22959: duty=91;
15'd22960: duty=102; 15'd22961: duty=105; 15'd22962: duty=112; 15'd22963: duty=107; 15'd22964: duty=107; 15'd22965: duty=107; 15'd22966: duty=100; 15'd22967: duty=107;
15'd22968: duty=110; 15'd22969: duty=116; 15'd22970: duty=106; 15'd22971: duty=112; 15'd22972: duty=107; 15'd22973: duty=114; 15'd22974: duty=126; 15'd22975: duty=111;
15'd22976: duty=115; 15'd22977: duty=109; 15'd22978: duty=114; 15'd22979: duty=128; 15'd22980: duty=127; 15'd22981: duty=123; 15'd22982: duty=129; 15'd22983: duty=134;
15'd22984: duty=136; 15'd22985: duty=135; 15'd22986: duty=136; 15'd22987: duty=134; 15'd22988: duty=138; 15'd22989: duty=132; 15'd22990: duty=135; 15'd22991: duty=150;
15'd22992: duty=148; 15'd22993: duty=152; 15'd22994: duty=153; 15'd22995: duty=157; 15'd22996: duty=157; 15'd22997: duty=157; 15'd22998: duty=145; 15'd22999: duty=143;
15'd23000: duty=141; 15'd23001: duty=148; 15'd23002: duty=154; 15'd23003: duty=148; 15'd23004: duty=156; 15'd23005: duty=152; 15'd23006: duty=157; 15'd23007: duty=160;
15'd23008: duty=166; 15'd23009: duty=165; 15'd23010: duty=159; 15'd23011: duty=157; 15'd23012: duty=163; 15'd23013: duty=153; 15'd23014: duty=151; 15'd23015: duty=150;
15'd23016: duty=139; 15'd23017: duty=142; 15'd23018: duty=138; 15'd23019: duty=156; 15'd23020: duty=139; 15'd23021: duty=136; 15'd23022: duty=140; 15'd23023: duty=142;
15'd23024: duty=137; 15'd23025: duty=139; 15'd23026: duty=135; 15'd23027: duty=126; 15'd23028: duty=122; 15'd23029: duty=108; 15'd23030: duty=110; 15'd23031: duty=103;
15'd23032: duty=101; 15'd23033: duty=107; 15'd23034: duty=97; 15'd23035: duty=102; 15'd23036: duty=110; 15'd23037: duty=95; 15'd23038: duty=115; 15'd23039: duty=107;
15'd23040: duty=107; 15'd23041: duty=107; 15'd23042: duty=99; 15'd23043: duty=101; 15'd23044: duty=98; 15'd23045: duty=93; 15'd23046: duty=90; 15'd23047: duty=96;
15'd23048: duty=99; 15'd23049: duty=104; 15'd23050: duty=102; 15'd23051: duty=110; 15'd23052: duty=122; 15'd23053: duty=122; 15'd23054: duty=118; 15'd23055: duty=124;
15'd23056: duty=122; 15'd23057: duty=125; 15'd23058: duty=133; 15'd23059: duty=125; 15'd23060: duty=133; 15'd23061: duty=136; 15'd23062: duty=133; 15'd23063: duty=134;
15'd23064: duty=142; 15'd23065: duty=145; 15'd23066: duty=146; 15'd23067: duty=134; 15'd23068: duty=132; 15'd23069: duty=142; 15'd23070: duty=146; 15'd23071: duty=160;
15'd23072: duty=151; 15'd23073: duty=154; 15'd23074: duty=161; 15'd23075: duty=163; 15'd23076: duty=163; 15'd23077: duty=162; 15'd23078: duty=172; 15'd23079: duty=174;
15'd23080: duty=159; 15'd23081: duty=158; 15'd23082: duty=146; 15'd23083: duty=138; 15'd23084: duty=140; 15'd23085: duty=135; 15'd23086: duty=140; 15'd23087: duty=152;
15'd23088: duty=151; 15'd23089: duty=158; 15'd23090: duty=163; 15'd23091: duty=155; 15'd23092: duty=152; 15'd23093: duty=142; 15'd23094: duty=135; 15'd23095: duty=132;
15'd23096: duty=134; 15'd23097: duty=132; 15'd23098: duty=134; 15'd23099: duty=123; 15'd23100: duty=123; 15'd23101: duty=125; 15'd23102: duty=123; 15'd23103: duty=121;
15'd23104: duty=123; 15'd23105: duty=120; 15'd23106: duty=117; 15'd23107: duty=115; 15'd23108: duty=107; 15'd23109: duty=117; 15'd23110: duty=120; 15'd23111: duty=103;
15'd23112: duty=97; 15'd23113: duty=100; 15'd23114: duty=106; 15'd23115: duty=111; 15'd23116: duty=113; 15'd23117: duty=112; 15'd23118: duty=104; 15'd23119: duty=93;
15'd23120: duty=93; 15'd23121: duty=96; 15'd23122: duty=100; 15'd23123: duty=96; 15'd23124: duty=91; 15'd23125: duty=106; 15'd23126: duty=105; 15'd23127: duty=115;
15'd23128: duty=124; 15'd23129: duty=119; 15'd23130: duty=128; 15'd23131: duty=128; 15'd23132: duty=122; 15'd23133: duty=121; 15'd23134: duty=113; 15'd23135: duty=118;
15'd23136: duty=116; 15'd23137: duty=116; 15'd23138: duty=123; 15'd23139: duty=118; 15'd23140: duty=124; 15'd23141: duty=134; 15'd23142: duty=139; 15'd23143: duty=146;
15'd23144: duty=151; 15'd23145: duty=160; 15'd23146: duty=170; 15'd23147: duty=182; 15'd23148: duty=173; 15'd23149: duty=181; 15'd23150: duty=178; 15'd23151: duty=175;
15'd23152: duty=178; 15'd23153: duty=169; 15'd23154: duty=170; 15'd23155: duty=159; 15'd23156: duty=166; 15'd23157: duty=154; 15'd23158: duty=156; 15'd23159: duty=161;
15'd23160: duty=151; 15'd23161: duty=154; 15'd23162: duty=153; 15'd23163: duty=152; 15'd23164: duty=165; 15'd23165: duty=157; 15'd23166: duty=150; 15'd23167: duty=149;
15'd23168: duty=139; 15'd23169: duty=137; 15'd23170: duty=139; 15'd23171: duty=135; 15'd23172: duty=142; 15'd23173: duty=139; 15'd23174: duty=126; 15'd23175: duty=125;
15'd23176: duty=130; 15'd23177: duty=132; 15'd23178: duty=119; 15'd23179: duty=108; 15'd23180: duty=103; 15'd23181: duty=116; 15'd23182: duty=116; 15'd23183: duty=102;
15'd23184: duty=101; 15'd23185: duty=103; 15'd23186: duty=104; 15'd23187: duty=98; 15'd23188: duty=83; 15'd23189: duty=98; 15'd23190: duty=92; 15'd23191: duty=88;
15'd23192: duty=96; 15'd23193: duty=101; 15'd23194: duty=107; 15'd23195: duty=92; 15'd23196: duty=103; 15'd23197: duty=98; 15'd23198: duty=90; 15'd23199: duty=89;
15'd23200: duty=95; 15'd23201: duty=98; 15'd23202: duty=102; 15'd23203: duty=112; 15'd23204: duty=98; 15'd23205: duty=119; 15'd23206: duty=122; 15'd23207: duty=116;
15'd23208: duty=127; 15'd23209: duty=123; 15'd23210: duty=131; 15'd23211: duty=124; 15'd23212: duty=127; 15'd23213: duty=134; 15'd23214: duty=139; 15'd23215: duty=139;
15'd23216: duty=140; 15'd23217: duty=149; 15'd23218: duty=149; 15'd23219: duty=156; 15'd23220: duty=157; 15'd23221: duty=157; 15'd23222: duty=159; 15'd23223: duty=154;
15'd23224: duty=156; 15'd23225: duty=161; 15'd23226: duty=163; 15'd23227: duty=156; 15'd23228: duty=154; 15'd23229: duty=159; 15'd23230: duty=165; 15'd23231: duty=165;
15'd23232: duty=161; 15'd23233: duty=165; 15'd23234: duty=153; 15'd23235: duty=158; 15'd23236: duty=162; 15'd23237: duty=162; 15'd23238: duty=159; 15'd23239: duty=157;
15'd23240: duty=148; 15'd23241: duty=149; 15'd23242: duty=156; 15'd23243: duty=152; 15'd23244: duty=152; 15'd23245: duty=139; 15'd23246: duty=142; 15'd23247: duty=145;
15'd23248: duty=142; 15'd23249: duty=139; 15'd23250: duty=132; 15'd23251: duty=125; 15'd23252: duty=129; 15'd23253: duty=135; 15'd23254: duty=125; 15'd23255: duty=126;
15'd23256: duty=123; 15'd23257: duty=112; 15'd23258: duty=108; 15'd23259: duty=101; 15'd23260: duty=105; 15'd23261: duty=106; 15'd23262: duty=110; 15'd23263: duty=114;
15'd23264: duty=109; 15'd23265: duty=102; 15'd23266: duty=97; 15'd23267: duty=98; 15'd23268: duty=105; 15'd23269: duty=98; 15'd23270: duty=100; 15'd23271: duty=103;
15'd23272: duty=111; 15'd23273: duty=111; 15'd23274: duty=106; 15'd23275: duty=108; 15'd23276: duty=97; 15'd23277: duty=91; 15'd23278: duty=89; 15'd23279: duty=95;
15'd23280: duty=102; 15'd23281: duty=112; 15'd23282: duty=107; 15'd23283: duty=112; 15'd23284: duty=116; 15'd23285: duty=118; 15'd23286: duty=126; 15'd23287: duty=126;
15'd23288: duty=125; 15'd23289: duty=132; 15'd23290: duty=131; 15'd23291: duty=124; 15'd23292: duty=131; 15'd23293: duty=126; 15'd23294: duty=127; 15'd23295: duty=128;
15'd23296: duty=132; 15'd23297: duty=142; 15'd23298: duty=151; 15'd23299: duty=143; 15'd23300: duty=148; 15'd23301: duty=148; 15'd23302: duty=148; 15'd23303: duty=165;
15'd23304: duty=162; 15'd23305: duty=154; 15'd23306: duty=145; 15'd23307: duty=153; 15'd23308: duty=163; 15'd23309: duty=171; 15'd23310: duty=162; 15'd23311: duty=160;
15'd23312: duty=164; 15'd23313: duty=165; 15'd23314: duty=168; 15'd23315: duty=171; 15'd23316: duty=171; 15'd23317: duty=162; 15'd23318: duty=160; 15'd23319: duty=166;
15'd23320: duty=166; 15'd23321: duty=153; 15'd23322: duty=158; 15'd23323: duty=148; 15'd23324: duty=142; 15'd23325: duty=150; 15'd23326: duty=148; 15'd23327: duty=150;
15'd23328: duty=137; 15'd23329: duty=136; 15'd23330: duty=139; 15'd23331: duty=126; 15'd23332: duty=128; 15'd23333: duty=124; 15'd23334: duty=124; 15'd23335: duty=115;
15'd23336: duty=105; 15'd23337: duty=102; 15'd23338: duty=99; 15'd23339: duty=98; 15'd23340: duty=108; 15'd23341: duty=112; 15'd23342: duty=107; 15'd23343: duty=97;
15'd23344: duty=103; 15'd23345: duty=109; 15'd23346: duty=102; 15'd23347: duty=94; 15'd23348: duty=88; 15'd23349: duty=97; 15'd23350: duty=94; 15'd23351: duty=100;
15'd23352: duty=94; 15'd23353: duty=95; 15'd23354: duty=97; 15'd23355: duty=106; 15'd23356: duty=115; 15'd23357: duty=106; 15'd23358: duty=100; 15'd23359: duty=112;
15'd23360: duty=117; 15'd23361: duty=117; 15'd23362: duty=120; 15'd23363: duty=119; 15'd23364: duty=120; 15'd23365: duty=119; 15'd23366: duty=126; 15'd23367: duty=122;
15'd23368: duty=130; 15'd23369: duty=138; 15'd23370: duty=140; 15'd23371: duty=141; 15'd23372: duty=141; 15'd23373: duty=130; 15'd23374: duty=132; 15'd23375: duty=143;
15'd23376: duty=141; 15'd23377: duty=144; 15'd23378: duty=146; 15'd23379: duty=142; 15'd23380: duty=149; 15'd23381: duty=159; 15'd23382: duty=160; 15'd23383: duty=167;
15'd23384: duty=165; 15'd23385: duty=171; 15'd23386: duty=174; 15'd23387: duty=167; 15'd23388: duty=160; 15'd23389: duty=161; 15'd23390: duty=159; 15'd23391: duty=157;
15'd23392: duty=155; 15'd23393: duty=154; 15'd23394: duty=168; 15'd23395: duty=163; 15'd23396: duty=164; 15'd23397: duty=167; 15'd23398: duty=159; 15'd23399: duty=161;
15'd23400: duty=153; 15'd23401: duty=148; 15'd23402: duty=139; 15'd23403: duty=137; 15'd23404: duty=135; 15'd23405: duty=129; 15'd23406: duty=135; 15'd23407: duty=133;
15'd23408: duty=132; 15'd23409: duty=125; 15'd23410: duty=123; 15'd23411: duty=132; 15'd23412: duty=132; 15'd23413: duty=125; 15'd23414: duty=117; 15'd23415: duty=114;
15'd23416: duty=119; 15'd23417: duty=111; 15'd23418: duty=114; 15'd23419: duty=100; 15'd23420: duty=100; 15'd23421: duty=96; 15'd23422: duty=89; 15'd23423: duty=108;
15'd23424: duty=95; 15'd23425: duty=96; 15'd23426: duty=94; 15'd23427: duty=96; 15'd23428: duty=104; 15'd23429: duty=106; 15'd23430: duty=105; 15'd23431: duty=108;
15'd23432: duty=106; 15'd23433: duty=104; 15'd23434: duty=100; 15'd23435: duty=100; 15'd23436: duty=106; 15'd23437: duty=113; 15'd23438: duty=104; 15'd23439: duty=105;
15'd23440: duty=112; 15'd23441: duty=113; 15'd23442: duty=122; 15'd23443: duty=114; 15'd23444: duty=110; 15'd23445: duty=120; 15'd23446: duty=128; 15'd23447: duty=129;
15'd23448: duty=134; 15'd23449: duty=139; 15'd23450: duty=133; 15'd23451: duty=136; 15'd23452: duty=147; 15'd23453: duty=153; 15'd23454: duty=158; 15'd23455: duty=156;
15'd23456: duty=158; 15'd23457: duty=162; 15'd23458: duty=154; 15'd23459: duty=149; 15'd23460: duty=159; 15'd23461: duty=163; 15'd23462: duty=159; 15'd23463: duty=155;
15'd23464: duty=164; 15'd23465: duty=165; 15'd23466: duty=175; 15'd23467: duty=174; 15'd23468: duty=176; 15'd23469: duty=171; 15'd23470: duty=175; 15'd23471: duty=172;
15'd23472: duty=167; 15'd23473: duty=174; 15'd23474: duty=166; 15'd23475: duty=166; 15'd23476: duty=158; 15'd23477: duty=146; 15'd23478: duty=152; 15'd23479: duty=151;
15'd23480: duty=138; 15'd23481: duty=146; 15'd23482: duty=133; 15'd23483: duty=138; 15'd23484: duty=135; 15'd23485: duty=132; 15'd23486: duty=123; 15'd23487: duty=123;
15'd23488: duty=109; 15'd23489: duty=109; 15'd23490: duty=122; 15'd23491: duty=113; 15'd23492: duty=106; 15'd23493: duty=102; 15'd23494: duty=106; 15'd23495: duty=88;
15'd23496: duty=86; 15'd23497: duty=88; 15'd23498: duty=106; 15'd23499: duty=97; 15'd23500: duty=97; 15'd23501: duty=93; 15'd23502: duty=86; 15'd23503: duty=92;
15'd23504: duty=88; 15'd23505: duty=110; 15'd23506: duty=109; 15'd23507: duty=93; 15'd23508: duty=92; 15'd23509: duty=90; 15'd23510: duty=92; 15'd23511: duty=101;
15'd23512: duty=98; 15'd23513: duty=93; 15'd23514: duty=101; 15'd23515: duty=102; 15'd23516: duty=105; 15'd23517: duty=110; 15'd23518: duty=110; 15'd23519: duty=116;
15'd23520: duty=116; 15'd23521: duty=119; 15'd23522: duty=125; 15'd23523: duty=130; 15'd23524: duty=131; 15'd23525: duty=130; 15'd23526: duty=134; 15'd23527: duty=139;
15'd23528: duty=136; 15'd23529: duty=145; 15'd23530: duty=155; 15'd23531: duty=159; 15'd23532: duty=154; 15'd23533: duty=150; 15'd23534: duty=163; 15'd23535: duty=168;
15'd23536: duty=180; 15'd23537: duty=185; 15'd23538: duty=175; 15'd23539: duty=173; 15'd23540: duty=166; 15'd23541: duty=167; 15'd23542: duty=171; 15'd23543: duty=168;
15'd23544: duty=166; 15'd23545: duty=164; 15'd23546: duty=165; 15'd23547: duty=164; 15'd23548: duty=168; 15'd23549: duty=170; 15'd23550: duty=168; 15'd23551: duty=165;
15'd23552: duty=168; 15'd23553: duty=156; 15'd23554: duty=157; 15'd23555: duty=160; 15'd23556: duty=159; 15'd23557: duty=146; 15'd23558: duty=139; 15'd23559: duty=134;
15'd23560: duty=133; 15'd23561: duty=132; 15'd23562: duty=128; 15'd23563: duty=132; 15'd23564: duty=118; 15'd23565: duty=116; 15'd23566: duty=118; 15'd23567: duty=119;
15'd23568: duty=124; 15'd23569: duty=116; 15'd23570: duty=104; 15'd23571: duty=113; 15'd23572: duty=94; 15'd23573: duty=105; 15'd23574: duty=120; 15'd23575: duty=105;
15'd23576: duty=103; 15'd23577: duty=91; 15'd23578: duty=100; 15'd23579: duty=90; 15'd23580: duty=91; 15'd23581: duty=88; 15'd23582: duty=92; 15'd23583: duty=90;
15'd23584: duty=75; 15'd23585: duty=102; 15'd23586: duty=95; 15'd23587: duty=96; 15'd23588: duty=104; 15'd23589: duty=102; 15'd23590: duty=107; 15'd23591: duty=110;
15'd23592: duty=113; 15'd23593: duty=114; 15'd23594: duty=115; 15'd23595: duty=105; 15'd23596: duty=107; 15'd23597: duty=116; 15'd23598: duty=119; 15'd23599: duty=119;
15'd23600: duty=107; 15'd23601: duty=115; 15'd23602: duty=121; 15'd23603: duty=124; 15'd23604: duty=133; 15'd23605: duty=129; 15'd23606: duty=136; 15'd23607: duty=143;
15'd23608: duty=143; 15'd23609: duty=151; 15'd23610: duty=162; 15'd23611: duty=166; 15'd23612: duty=165; 15'd23613: duty=157; 15'd23614: duty=156; 15'd23615: duty=152;
15'd23616: duty=159; 15'd23617: duty=154; 15'd23618: duty=153; 15'd23619: duty=149; 15'd23620: duty=156; 15'd23621: duty=159; 15'd23622: duty=159; 15'd23623: duty=174;
15'd23624: duty=167; 15'd23625: duty=183; 15'd23626: duty=173; 15'd23627: duty=162; 15'd23628: duty=173; 15'd23629: duty=166; 15'd23630: duty=161; 15'd23631: duty=159;
15'd23632: duty=151; 15'd23633: duty=149; 15'd23634: duty=156; 15'd23635: duty=157; 15'd23636: duty=149; 15'd23637: duty=148; 15'd23638: duty=141; 15'd23639: duty=140;
15'd23640: duty=135; 15'd23641: duty=125; 15'd23642: duty=126; 15'd23643: duty=135; 15'd23644: duty=133; 15'd23645: duty=125; 15'd23646: duty=123; 15'd23647: duty=119;
15'd23648: duty=127; 15'd23649: duty=119; 15'd23650: duty=113; 15'd23651: duty=107; 15'd23652: duty=93; 15'd23653: duty=93; 15'd23654: duty=93; 15'd23655: duty=96;
15'd23656: duty=89; 15'd23657: duty=86; 15'd23658: duty=91; 15'd23659: duty=87; 15'd23660: duty=104; 15'd23661: duty=102; 15'd23662: duty=106; 15'd23663: duty=104;
15'd23664: duty=94; 15'd23665: duty=87; 15'd23666: duty=93; 15'd23667: duty=111; 15'd23668: duty=112; 15'd23669: duty=110; 15'd23670: duty=107; 15'd23671: duty=113;
15'd23672: duty=115; 15'd23673: duty=107; 15'd23674: duty=109; 15'd23675: duty=115; 15'd23676: duty=115; 15'd23677: duty=121; 15'd23678: duty=121; 15'd23679: duty=134;
15'd23680: duty=136; 15'd23681: duty=124; 15'd23682: duty=128; 15'd23683: duty=137; 15'd23684: duty=148; 15'd23685: duty=154; 15'd23686: duty=153; 15'd23687: duty=160;
15'd23688: duty=157; 15'd23689: duty=162; 15'd23690: duty=151; 15'd23691: duty=150; 15'd23692: duty=155; 15'd23693: duty=156; 15'd23694: duty=152; 15'd23695: duty=153;
15'd23696: duty=165; 15'd23697: duty=155; 15'd23698: duty=160; 15'd23699: duty=164; 15'd23700: duty=158; 15'd23701: duty=161; 15'd23702: duty=165; 15'd23703: duty=162;
15'd23704: duty=166; 15'd23705: duty=168; 15'd23706: duty=160; 15'd23707: duty=147; 15'd23708: duty=146; 15'd23709: duty=139; 15'd23710: duty=138; 15'd23711: duty=131;
15'd23712: duty=135; 15'd23713: duty=138; 15'd23714: duty=134; 15'd23715: duty=141; 15'd23716: duty=134; 15'd23717: duty=133; 15'd23718: duty=132; 15'd23719: duty=133;
15'd23720: duty=132; 15'd23721: duty=134; 15'd23722: duty=127; 15'd23723: duty=120; 15'd23724: duty=117; 15'd23725: duty=115; 15'd23726: duty=118; 15'd23727: duty=113;
15'd23728: duty=113; 15'd23729: duty=107; 15'd23730: duty=102; 15'd23731: duty=99; 15'd23732: duty=107; 15'd23733: duty=110; 15'd23734: duty=99; 15'd23735: duty=102;
15'd23736: duty=107; 15'd23737: duty=109; 15'd23738: duty=105; 15'd23739: duty=112; 15'd23740: duty=105; 15'd23741: duty=107; 15'd23742: duty=113; 15'd23743: duty=114;
15'd23744: duty=118; 15'd23745: duty=115; 15'd23746: duty=107; 15'd23747: duty=108; 15'd23748: duty=115; 15'd23749: duty=108; 15'd23750: duty=108; 15'd23751: duty=118;
15'd23752: duty=121; 15'd23753: duty=116; 15'd23754: duty=124; 15'd23755: duty=118; 15'd23756: duty=119; 15'd23757: duty=121; 15'd23758: duty=127; 15'd23759: duty=140;
15'd23760: duty=141; 15'd23761: duty=140; 15'd23762: duty=141; 15'd23763: duty=149; 15'd23764: duty=147; 15'd23765: duty=154; 15'd23766: duty=150; 15'd23767: duty=141;
15'd23768: duty=147; 15'd23769: duty=149; 15'd23770: duty=156; 15'd23771: duty=147; 15'd23772: duty=159; 15'd23773: duty=163; 15'd23774: duty=158; 15'd23775: duty=162;
15'd23776: duty=165; 15'd23777: duty=169; 15'd23778: duty=157; 15'd23779: duty=160; 15'd23780: duty=162; 15'd23781: duty=162; 15'd23782: duty=157; 15'd23783: duty=151;
15'd23784: duty=148; 15'd23785: duty=146; 15'd23786: duty=142; 15'd23787: duty=151; 15'd23788: duty=153; 15'd23789: duty=139; 15'd23790: duty=141; 15'd23791: duty=145;
15'd23792: duty=128; 15'd23793: duty=132; 15'd23794: duty=135; 15'd23795: duty=131; 15'd23796: duty=131; 15'd23797: duty=115; 15'd23798: duty=121; 15'd23799: duty=116;
15'd23800: duty=110; 15'd23801: duty=107; 15'd23802: duty=108; 15'd23803: duty=113; 15'd23804: duty=108; 15'd23805: duty=115; 15'd23806: duty=122; 15'd23807: duty=116;
15'd23808: duty=107; 15'd23809: duty=102; 15'd23810: duty=102; 15'd23811: duty=113; 15'd23812: duty=113; 15'd23813: duty=109; 15'd23814: duty=121; 15'd23815: duty=110;
15'd23816: duty=104; 15'd23817: duty=107; 15'd23818: duty=110; 15'd23819: duty=112; 15'd23820: duty=119; 15'd23821: duty=119; 15'd23822: duty=107; 15'd23823: duty=103;
15'd23824: duty=100; 15'd23825: duty=104; 15'd23826: duty=116; 15'd23827: duty=123; 15'd23828: duty=121; 15'd23829: duty=127; 15'd23830: duty=128; 15'd23831: duty=133;
15'd23832: duty=135; 15'd23833: duty=137; 15'd23834: duty=129; 15'd23835: duty=130; 15'd23836: duty=135; 15'd23837: duty=142; 15'd23838: duty=149; 15'd23839: duty=144;
15'd23840: duty=149; 15'd23841: duty=146; 15'd23842: duty=150; 15'd23843: duty=158; 15'd23844: duty=161; 15'd23845: duty=159; 15'd23846: duty=154; 15'd23847: duty=150;
15'd23848: duty=154; 15'd23849: duty=150; 15'd23850: duty=158; 15'd23851: duty=155; 15'd23852: duty=154; 15'd23853: duty=158; 15'd23854: duty=164; 15'd23855: duty=161;
15'd23856: duty=160; 15'd23857: duty=164; 15'd23858: duty=145; 15'd23859: duty=153; 15'd23860: duty=152; 15'd23861: duty=153; 15'd23862: duty=143; 15'd23863: duty=138;
15'd23864: duty=138; 15'd23865: duty=139; 15'd23866: duty=141; 15'd23867: duty=136; 15'd23868: duty=129; 15'd23869: duty=121; 15'd23870: duty=128; 15'd23871: duty=131;
15'd23872: duty=127; 15'd23873: duty=126; 15'd23874: duty=127; 15'd23875: duty=119; 15'd23876: duty=116; 15'd23877: duty=110; 15'd23878: duty=118; 15'd23879: duty=115;
15'd23880: duty=113; 15'd23881: duty=113; 15'd23882: duty=113; 15'd23883: duty=116; 15'd23884: duty=118; 15'd23885: duty=115; 15'd23886: duty=104; 15'd23887: duty=101;
15'd23888: duty=109; 15'd23889: duty=104; 15'd23890: duty=94; 15'd23891: duty=105; 15'd23892: duty=99; 15'd23893: duty=104; 15'd23894: duty=112; 15'd23895: duty=109;
15'd23896: duty=96; 15'd23897: duty=98; 15'd23898: duty=101; 15'd23899: duty=102; 15'd23900: duty=107; 15'd23901: duty=112; 15'd23902: duty=117; 15'd23903: duty=114;
15'd23904: duty=114; 15'd23905: duty=118; 15'd23906: duty=125; 15'd23907: duty=118; 15'd23908: duty=119; 15'd23909: duty=121; 15'd23910: duty=128; 15'd23911: duty=142;
15'd23912: duty=138; 15'd23913: duty=141; 15'd23914: duty=152; 15'd23915: duty=154; 15'd23916: duty=158; 15'd23917: duty=164; 15'd23918: duty=155; 15'd23919: duty=150;
15'd23920: duty=142; 15'd23921: duty=144; 15'd23922: duty=148; 15'd23923: duty=145; 15'd23924: duty=150; 15'd23925: duty=154; 15'd23926: duty=162; 15'd23927: duty=160;
15'd23928: duty=165; 15'd23929: duty=160; 15'd23930: duty=158; 15'd23931: duty=155; 15'd23932: duty=155; 15'd23933: duty=166; 15'd23934: duty=171; 15'd23935: duty=165;
15'd23936: duty=156; 15'd23937: duty=149; 15'd23938: duty=141; 15'd23939: duty=141; 15'd23940: duty=141; 15'd23941: duty=138; 15'd23942: duty=140; 15'd23943: duty=149;
15'd23944: duty=142; 15'd23945: duty=140; 15'd23946: duty=135; 15'd23947: duty=130; 15'd23948: duty=136; 15'd23949: duty=137; 15'd23950: duty=126; 15'd23951: duty=128;
15'd23952: duty=118; 15'd23953: duty=113; 15'd23954: duty=106; 15'd23955: duty=99; 15'd23956: duty=108; 15'd23957: duty=99; 15'd23958: duty=104; 15'd23959: duty=110;
15'd23960: duty=112; 15'd23961: duty=104; 15'd23962: duty=99; 15'd23963: duty=101; 15'd23964: duty=104; 15'd23965: duty=104; 15'd23966: duty=99; 15'd23967: duty=99;
15'd23968: duty=108; 15'd23969: duty=108; 15'd23970: duty=111; 15'd23971: duty=109; 15'd23972: duty=112; 15'd23973: duty=115; 15'd23974: duty=116; 15'd23975: duty=117;
15'd23976: duty=116; 15'd23977: duty=130; 15'd23978: duty=135; 15'd23979: duty=131; 15'd23980: duty=125; 15'd23981: duty=126; 15'd23982: duty=125; 15'd23983: duty=135;
15'd23984: duty=138; 15'd23985: duty=136; 15'd23986: duty=131; 15'd23987: duty=131; 15'd23988: duty=138; 15'd23989: duty=148; 15'd23990: duty=141; 15'd23991: duty=130;
15'd23992: duty=140; 15'd23993: duty=145; 15'd23994: duty=151; 15'd23995: duty=154; 15'd23996: duty=158; 15'd23997: duty=157; 15'd23998: duty=157; 15'd23999: duty=142;
15'd24000: duty=139; 15'd24001: duty=147; 15'd24002: duty=148; 15'd24003: duty=149; 15'd24004: duty=153; 15'd24005: duty=151; 15'd24006: duty=150; 15'd24007: duty=146;
15'd24008: duty=141; 15'd24009: duty=137; 15'd24010: duty=128; 15'd24011: duty=132; 15'd24012: duty=131; 15'd24013: duty=143; 15'd24014: duty=134; 15'd24015: duty=134;
15'd24016: duty=131; 15'd24017: duty=132; 15'd24018: duty=133; 15'd24019: duty=122; 15'd24020: duty=128; 15'd24021: duty=122; 15'd24022: duty=136; 15'd24023: duty=131;
15'd24024: duty=122; 15'd24025: duty=127; 15'd24026: duty=126; 15'd24027: duty=116; 15'd24028: duty=127; 15'd24029: duty=129; 15'd24030: duty=118; 15'd24031: duty=111;
15'd24032: duty=108; 15'd24033: duty=122; 15'd24034: duty=121; 15'd24035: duty=124; 15'd24036: duty=121; 15'd24037: duty=127; 15'd24038: duty=131; 15'd24039: duty=127;
15'd24040: duty=125; 15'd24041: duty=110; 15'd24042: duty=107; 15'd24043: duty=112; 15'd24044: duty=117; 15'd24045: duty=115; 15'd24046: duty=111; 15'd24047: duty=128;
15'd24048: duty=124; 15'd24049: duty=128; 15'd24050: duty=122; 15'd24051: duty=130; 15'd24052: duty=132; 15'd24053: duty=136; 15'd24054: duty=145; 15'd24055: duty=139;
15'd24056: duty=142; 15'd24057: duty=136; 15'd24058: duty=137; 15'd24059: duty=120; 15'd24060: duty=117; 15'd24061: duty=118; 15'd24062: duty=123; 15'd24063: duty=124;
15'd24064: duty=128; 15'd24065: duty=133; 15'd24066: duty=140; 15'd24067: duty=145; 15'd24068: duty=142; 15'd24069: duty=141; 15'd24070: duty=140; 15'd24071: duty=142;
15'd24072: duty=139; 15'd24073: duty=134; 15'd24074: duty=142; 15'd24075: duty=139; 15'd24076: duty=139; 15'd24077: duty=136; 15'd24078: duty=142; 15'd24079: duty=146;
15'd24080: duty=142; 15'd24081: duty=150; 15'd24082: duty=144; 15'd24083: duty=148; 15'd24084: duty=149; 15'd24085: duty=152; 15'd24086: duty=144; 15'd24087: duty=145;
15'd24088: duty=144; 15'd24089: duty=134; 15'd24090: duty=138; 15'd24091: duty=136; 15'd24092: duty=133; 15'd24093: duty=139; 15'd24094: duty=139; 15'd24095: duty=142;
15'd24096: duty=135; 15'd24097: duty=130; 15'd24098: duty=130; 15'd24099: duty=125; 15'd24100: duty=121; 15'd24101: duty=123; 15'd24102: duty=124; 15'd24103: duty=126;
15'd24104: duty=122; 15'd24105: duty=123; 15'd24106: duty=120; 15'd24107: duty=104; 15'd24108: duty=109; 15'd24109: duty=124; 15'd24110: duty=113; 15'd24111: duty=107;
15'd24112: duty=118; 15'd24113: duty=116; 15'd24114: duty=116; 15'd24115: duty=105; 15'd24116: duty=95; 15'd24117: duty=98; 15'd24118: duty=104; 15'd24119: duty=101;
15'd24120: duty=110; 15'd24121: duty=129; 15'd24122: duty=131; 15'd24123: duty=118; 15'd24124: duty=122; 15'd24125: duty=126; 15'd24126: duty=137; 15'd24127: duty=134;
15'd24128: duty=127; 15'd24129: duty=126; 15'd24130: duty=121; 15'd24131: duty=124; 15'd24132: duty=116; 15'd24133: duty=126; 15'd24134: duty=124; 15'd24135: duty=126;
15'd24136: duty=128; 15'd24137: duty=130; 15'd24138: duty=131; 15'd24139: duty=138; 15'd24140: duty=145; 15'd24141: duty=151; 15'd24142: duty=152; 15'd24143: duty=158;
15'd24144: duty=157; 15'd24145: duty=148; 15'd24146: duty=145; 15'd24147: duty=145; 15'd24148: duty=146; 15'd24149: duty=148; 15'd24150: duty=147; 15'd24151: duty=142;
15'd24152: duty=151; 15'd24153: duty=146; 15'd24154: duty=153; 15'd24155: duty=159; 15'd24156: duty=159; 15'd24157: duty=159; 15'd24158: duty=162; 15'd24159: duty=163;
15'd24160: duty=158; 15'd24161: duty=154; 15'd24162: duty=150; 15'd24163: duty=148; 15'd24164: duty=144; 15'd24165: duty=138; 15'd24166: duty=142; 15'd24167: duty=149;
15'd24168: duty=145; 15'd24169: duty=143; 15'd24170: duty=142; 15'd24171: duty=141; 15'd24172: duty=135; 15'd24173: duty=135; 15'd24174: duty=133; 15'd24175: duty=125;
15'd24176: duty=121; 15'd24177: duty=118; 15'd24178: duty=127; 15'd24179: duty=127; 15'd24180: duty=117; 15'd24181: duty=115; 15'd24182: duty=106; 15'd24183: duty=100;
15'd24184: duty=109; 15'd24185: duty=103; 15'd24186: duty=100; 15'd24187: duty=105; 15'd24188: duty=96; 15'd24189: duty=94; 15'd24190: duty=99; 15'd24191: duty=100;
15'd24192: duty=98; 15'd24193: duty=97; 15'd24194: duty=88; 15'd24195: duty=91; 15'd24196: duty=103; 15'd24197: duty=92; 15'd24198: duty=98; 15'd24199: duty=94;
15'd24200: duty=98; 15'd24201: duty=112; 15'd24202: duty=106; 15'd24203: duty=106; 15'd24204: duty=110; 15'd24205: duty=111; 15'd24206: duty=111; 15'd24207: duty=116;
15'd24208: duty=114; 15'd24209: duty=111; 15'd24210: duty=123; 15'd24211: duty=128; 15'd24212: duty=126; 15'd24213: duty=129; 15'd24214: duty=135; 15'd24215: duty=145;
15'd24216: duty=150; 15'd24217: duty=157; 15'd24218: duty=161; 15'd24219: duty=168; 15'd24220: duty=166; 15'd24221: duty=169; 15'd24222: duty=164; 15'd24223: duty=166;
15'd24224: duty=170; 15'd24225: duty=158; 15'd24226: duty=158; 15'd24227: duty=157; 15'd24228: duty=167; 15'd24229: duty=172; 15'd24230: duty=183; 15'd24231: duty=186;
15'd24232: duty=181; 15'd24233: duty=184; 15'd24234: duty=184; 15'd24235: duty=184; 15'd24236: duty=180; 15'd24237: duty=170; 15'd24238: duty=176; 15'd24239: duty=169;
15'd24240: duty=158; 15'd24241: duty=163; 15'd24242: duty=155; 15'd24243: duty=149; 15'd24244: duty=144; 15'd24245: duty=146; 15'd24246: duty=142; 15'd24247: duty=137;
15'd24248: duty=132; 15'd24249: duty=132; 15'd24250: duty=126; 15'd24251: duty=120; 15'd24252: duty=120; 15'd24253: duty=123; 15'd24254: duty=112; 15'd24255: duty=107;
15'd24256: duty=106; 15'd24257: duty=97; 15'd24258: duty=92; 15'd24259: duty=85; 15'd24260: duty=86; 15'd24261: duty=79; 15'd24262: duty=76; 15'd24263: duty=79;
15'd24264: duty=87; 15'd24265: duty=93; 15'd24266: duty=104; 15'd24267: duty=85; 15'd24268: duty=85; 15'd24269: duty=91; 15'd24270: duty=75; 15'd24271: duty=81;
15'd24272: duty=82; 15'd24273: duty=79; 15'd24274: duty=83; 15'd24275: duty=93; 15'd24276: duty=101; 15'd24277: duty=105; 15'd24278: duty=104; 15'd24279: duty=101;
15'd24280: duty=104; 15'd24281: duty=110; 15'd24282: duty=113; 15'd24283: duty=110; 15'd24284: duty=123; 15'd24285: duty=129; 15'd24286: duty=126; 15'd24287: duty=132;
15'd24288: duty=134; 15'd24289: duty=135; 15'd24290: duty=130; 15'd24291: duty=140; 15'd24292: duty=144; 15'd24293: duty=149; 15'd24294: duty=150; 15'd24295: duty=143;
15'd24296: duty=156; 15'd24297: duty=163; 15'd24298: duty=170; 15'd24299: duty=169; 15'd24300: duty=167; 15'd24301: duty=174; 15'd24302: duty=178; 15'd24303: duty=174;
15'd24304: duty=173; 15'd24305: duty=182; 15'd24306: duty=176; 15'd24307: duty=174; 15'd24308: duty=173; 15'd24309: duty=180; 15'd24310: duty=181; 15'd24311: duty=174;
15'd24312: duty=164; 15'd24313: duty=173; 15'd24314: duty=168; 15'd24315: duty=165; 15'd24316: duty=165; 15'd24317: duty=162; 15'd24318: duty=153; 15'd24319: duty=148;
15'd24320: duty=151; 15'd24321: duty=154; 15'd24322: duty=159; 15'd24323: duty=145; 15'd24324: duty=151; 15'd24325: duty=134; 15'd24326: duty=129; 15'd24327: duty=121;
15'd24328: duty=124; 15'd24329: duty=120; 15'd24330: duty=122; 15'd24331: duty=112; 15'd24332: duty=108; 15'd24333: duty=118; 15'd24334: duty=110; 15'd24335: duty=107;
15'd24336: duty=103; 15'd24337: duty=104; 15'd24338: duty=100; 15'd24339: duty=99; 15'd24340: duty=102; 15'd24341: duty=110; 15'd24342: duty=105; 15'd24343: duty=101;
15'd24344: duty=87; 15'd24345: duty=89; 15'd24346: duty=88; 15'd24347: duty=90; 15'd24348: duty=90; 15'd24349: duty=92; 15'd24350: duty=97; 15'd24351: duty=99;
15'd24352: duty=96; 15'd24353: duty=99; 15'd24354: duty=98; 15'd24355: duty=95; 15'd24356: duty=96; 15'd24357: duty=94; 15'd24358: duty=109; 15'd24359: duty=113;
15'd24360: duty=117; 15'd24361: duty=122; 15'd24362: duty=118; 15'd24363: duty=114; 15'd24364: duty=113; 15'd24365: duty=120; 15'd24366: duty=124; 15'd24367: duty=132;
15'd24368: duty=137; 15'd24369: duty=139; 15'd24370: duty=141; 15'd24371: duty=146; 15'd24372: duty=144; 15'd24373: duty=157; 15'd24374: duty=159; 15'd24375: duty=146;
15'd24376: duty=150; 15'd24377: duty=143; 15'd24378: duty=157; 15'd24379: duty=159; 15'd24380: duty=149; 15'd24381: duty=156; 15'd24382: duty=159; 15'd24383: duty=160;
15'd24384: duty=166; 15'd24385: duty=167; 15'd24386: duty=166; 15'd24387: duty=162; 15'd24388: duty=161; 15'd24389: duty=159; 15'd24390: duty=161; 15'd24391: duty=158;
15'd24392: duty=155; 15'd24393: duty=158; 15'd24394: duty=157; 15'd24395: duty=159; 15'd24396: duty=149; 15'd24397: duty=155; 15'd24398: duty=160; 15'd24399: duty=153;
15'd24400: duty=157; 15'd24401: duty=135; 15'd24402: duty=132; 15'd24403: duty=125; 15'd24404: duty=125; 15'd24405: duty=129; 15'd24406: duty=128; 15'd24407: duty=127;
15'd24408: duty=115; 15'd24409: duty=123; 15'd24410: duty=112; 15'd24411: duty=121; 15'd24412: duty=109; 15'd24413: duty=106; 15'd24414: duty=103; 15'd24415: duty=112;
15'd24416: duty=112; 15'd24417: duty=95; 15'd24418: duty=100; 15'd24419: duty=97; 15'd24420: duty=100; 15'd24421: duty=98; 15'd24422: duty=96; 15'd24423: duty=106;
15'd24424: duty=105; 15'd24425: duty=104; 15'd24426: duty=110; 15'd24427: duty=112; 15'd24428: duty=117; 15'd24429: duty=110; 15'd24430: duty=111; 15'd24431: duty=106;
15'd24432: duty=115; 15'd24433: duty=121; 15'd24434: duty=125; 15'd24435: duty=126; 15'd24436: duty=125; 15'd24437: duty=131; 15'd24438: duty=129; 15'd24439: duty=129;
15'd24440: duty=133; 15'd24441: duty=127; 15'd24442: duty=126; 15'd24443: duty=129; 15'd24444: duty=136; 15'd24445: duty=143; 15'd24446: duty=141; 15'd24447: duty=142;
15'd24448: duty=143; 15'd24449: duty=147; 15'd24450: duty=157; 15'd24451: duty=174; 15'd24452: duty=169; 15'd24453: duty=165; 15'd24454: duty=162; 15'd24455: duty=158;
15'd24456: duty=162; 15'd24457: duty=160; 15'd24458: duty=151; 15'd24459: duty=159; 15'd24460: duty=156; 15'd24461: duty=156; 15'd24462: duty=164; 15'd24463: duty=167;
15'd24464: duty=165; 15'd24465: duty=157; 15'd24466: duty=149; 15'd24467: duty=147; 15'd24468: duty=148; 15'd24469: duty=145; 15'd24470: duty=147; 15'd24471: duty=134;
15'd24472: duty=129; 15'd24473: duty=127; 15'd24474: duty=131; 15'd24475: duty=136; 15'd24476: duty=132; 15'd24477: duty=131; 15'd24478: duty=119; 15'd24479: duty=125;
15'd24480: duty=117; 15'd24481: duty=107; 15'd24482: duty=111; 15'd24483: duty=95; 15'd24484: duty=105; 15'd24485: duty=103; 15'd24486: duty=118; 15'd24487: duty=115;
15'd24488: duty=105; 15'd24489: duty=96; 15'd24490: duty=88; 15'd24491: duty=107; 15'd24492: duty=104; 15'd24493: duty=112; 15'd24494: duty=99; 15'd24495: duty=98;
15'd24496: duty=106; 15'd24497: duty=98; 15'd24498: duty=102; 15'd24499: duty=92; 15'd24500: duty=89; 15'd24501: duty=84; 15'd24502: duty=96; 15'd24503: duty=100;
15'd24504: duty=98; 15'd24505: duty=103; 15'd24506: duty=106; 15'd24507: duty=109; 15'd24508: duty=106; 15'd24509: duty=116; 15'd24510: duty=121; 15'd24511: duty=126;
15'd24512: duty=117; 15'd24513: duty=118; 15'd24514: duty=125; 15'd24515: duty=126; 15'd24516: duty=122; 15'd24517: duty=121; 15'd24518: duty=133; 15'd24519: duty=134;
15'd24520: duty=140; 15'd24521: duty=153; 15'd24522: duty=153; 15'd24523: duty=159; 15'd24524: duty=154; 15'd24525: duty=164; 15'd24526: duty=160; 15'd24527: duty=154;
15'd24528: duty=153; 15'd24529: duty=153; 15'd24530: duty=159; 15'd24531: duty=159; 15'd24532: duty=176; 15'd24533: duty=177; 15'd24534: duty=177; 15'd24535: duty=185;
15'd24536: duty=195; 15'd24537: duty=192; 15'd24538: duty=184; 15'd24539: duty=172; 15'd24540: duty=177; 15'd24541: duty=174; 15'd24542: duty=174; 15'd24543: duty=169;
15'd24544: duty=165; 15'd24545: duty=157; 15'd24546: duty=156; 15'd24547: duty=159; 15'd24548: duty=150; 15'd24549: duty=160; 15'd24550: duty=151; 15'd24551: duty=148;
15'd24552: duty=141; 15'd24553: duty=139; 15'd24554: duty=139; 15'd24555: duty=135; 15'd24556: duty=128; 15'd24557: duty=121; 15'd24558: duty=120; 15'd24559: duty=110;
15'd24560: duty=118; 15'd24561: duty=104; 15'd24562: duty=98; 15'd24563: duty=101; 15'd24564: duty=115; 15'd24565: duty=103; 15'd24566: duty=105; 15'd24567: duty=107;
15'd24568: duty=89; 15'd24569: duty=105; 15'd24570: duty=80; 15'd24571: duty=97; 15'd24572: duty=87; 15'd24573: duty=85; 15'd24574: duty=98; 15'd24575: duty=91;
15'd24576: duty=97; 15'd24577: duty=93; 15'd24578: duty=98; 15'd24579: duty=96; 15'd24580: duty=93; 15'd24581: duty=96; 15'd24582: duty=110; 15'd24583: duty=110;
15'd24584: duty=112; 15'd24585: duty=107; 15'd24586: duty=101; 15'd24587: duty=100; 15'd24588: duty=101; 15'd24589: duty=113; 15'd24590: duty=115; 15'd24591: duty=117;
15'd24592: duty=113; 15'd24593: duty=108; 15'd24594: duty=121; 15'd24595: duty=121; 15'd24596: duty=127; 15'd24597: duty=124; 15'd24598: duty=126; 15'd24599: duty=140;
15'd24600: duty=147; 15'd24601: duty=152; 15'd24602: duty=156; 15'd24603: duty=162; 15'd24604: duty=154; 15'd24605: duty=155; 15'd24606: duty=155; 15'd24607: duty=157;
15'd24608: duty=154; 15'd24609: duty=156; 15'd24610: duty=156; 15'd24611: duty=161; 15'd24612: duty=167; 15'd24613: duty=163; 15'd24614: duty=172; 15'd24615: duty=174;
15'd24616: duty=170; 15'd24617: duty=169; 15'd24618: duty=164; 15'd24619: duty=157; 15'd24620: duty=156; 15'd24621: duty=163; 15'd24622: duty=165; 15'd24623: duty=154;
15'd24624: duty=159; 15'd24625: duty=163; 15'd24626: duty=159; 15'd24627: duty=157; 15'd24628: duty=150; 15'd24629: duty=149; 15'd24630: duty=136; 15'd24631: duty=131;
15'd24632: duty=134; 15'd24633: duty=131; 15'd24634: duty=127; 15'd24635: duty=132; 15'd24636: duty=126; 15'd24637: duty=115; 15'd24638: duty=118; 15'd24639: duty=122;
15'd24640: duty=118; 15'd24641: duty=108; 15'd24642: duty=110; 15'd24643: duty=113; 15'd24644: duty=115; 15'd24645: duty=101; 15'd24646: duty=109; 15'd24647: duty=105;
15'd24648: duty=90; 15'd24649: duty=93; 15'd24650: duty=92; 15'd24651: duty=91; 15'd24652: duty=87; 15'd24653: duty=92; 15'd24654: duty=107; 15'd24655: duty=110;
15'd24656: duty=107; 15'd24657: duty=113; 15'd24658: duty=118; 15'd24659: duty=121; 15'd24660: duty=118; 15'd24661: duty=118; 15'd24662: duty=118; 15'd24663: duty=110;
15'd24664: duty=102; 15'd24665: duty=104; 15'd24666: duty=116; 15'd24667: duty=122; 15'd24668: duty=122; 15'd24669: duty=121; 15'd24670: duty=121; 15'd24671: duty=128;
15'd24672: duty=137; 15'd24673: duty=142; 15'd24674: duty=145; 15'd24675: duty=144; 15'd24676: duty=146; 15'd24677: duty=145; 15'd24678: duty=137; 15'd24679: duty=145;
15'd24680: duty=140; 15'd24681: duty=145; 15'd24682: duty=151; 15'd24683: duty=150; 15'd24684: duty=146; 15'd24685: duty=145; 15'd24686: duty=146; 15'd24687: duty=151;
15'd24688: duty=160; 15'd24689: duty=156; 15'd24690: duty=162; 15'd24691: duty=154; 15'd24692: duty=156; 15'd24693: duty=160; 15'd24694: duty=154; 15'd24695: duty=158;
15'd24696: duty=148; 15'd24697: duty=145; 15'd24698: duty=144; 15'd24699: duty=140; 15'd24700: duty=154; 15'd24701: duty=151; 15'd24702: duty=153; 15'd24703: duty=149;
15'd24704: duty=135; 15'd24705: duty=136; 15'd24706: duty=135; 15'd24707: duty=137; 15'd24708: duty=134; 15'd24709: duty=140; 15'd24710: duty=127; 15'd24711: duty=122;
15'd24712: duty=117; 15'd24713: duty=111; 15'd24714: duty=123; 15'd24715: duty=108; 15'd24716: duty=109; 15'd24717: duty=105; 15'd24718: duty=104; 15'd24719: duty=119;
15'd24720: duty=114; 15'd24721: duty=105; 15'd24722: duty=103; 15'd24723: duty=102; 15'd24724: duty=100; 15'd24725: duty=113; 15'd24726: duty=120; 15'd24727: duty=114;
15'd24728: duty=119; 15'd24729: duty=117; 15'd24730: duty=111; 15'd24731: duty=114; 15'd24732: duty=117; 15'd24733: duty=119; 15'd24734: duty=106; 15'd24735: duty=114;
15'd24736: duty=118; 15'd24737: duty=111; 15'd24738: duty=110; 15'd24739: duty=110; 15'd24740: duty=120; 15'd24741: duty=125; 15'd24742: duty=131; 15'd24743: duty=131;
15'd24744: duty=131; 15'd24745: duty=132; 15'd24746: duty=136; 15'd24747: duty=136; 15'd24748: duty=126; 15'd24749: duty=125; 15'd24750: duty=136; 15'd24751: duty=149;
15'd24752: duty=145; 15'd24753: duty=145; 15'd24754: duty=150; 15'd24755: duty=151; 15'd24756: duty=157; 15'd24757: duty=151; 15'd24758: duty=149; 15'd24759: duty=147;
15'd24760: duty=148; 15'd24761: duty=156; 15'd24762: duty=163; 15'd24763: duty=168; 15'd24764: duty=160; 15'd24765: duty=159; 15'd24766: duty=160; 15'd24767: duty=157;
15'd24768: duty=160; 15'd24769: duty=160; 15'd24770: duty=162; 15'd24771: duty=159; 15'd24772: duty=151; 15'd24773: duty=143; 15'd24774: duty=142; 15'd24775: duty=137;
15'd24776: duty=137; 15'd24777: duty=136; 15'd24778: duty=139; 15'd24779: duty=136; 15'd24780: duty=134; 15'd24781: duty=134; 15'd24782: duty=136; 15'd24783: duty=130;
15'd24784: duty=115; 15'd24785: duty=116; 15'd24786: duty=115; 15'd24787: duty=121; 15'd24788: duty=116; 15'd24789: duty=113; 15'd24790: duty=113; 15'd24791: duty=107;
15'd24792: duty=99; 15'd24793: duty=112; 15'd24794: duty=115; 15'd24795: duty=115; 15'd24796: duty=122; 15'd24797: duty=112; 15'd24798: duty=118; 15'd24799: duty=116;
15'd24800: duty=102; 15'd24801: duty=106; 15'd24802: duty=107; 15'd24803: duty=103; 15'd24804: duty=97; 15'd24805: duty=95; 15'd24806: duty=100; 15'd24807: duty=107;
15'd24808: duty=111; 15'd24809: duty=115; 15'd24810: duty=116; 15'd24811: duty=113; 15'd24812: duty=116; 15'd24813: duty=113; 15'd24814: duty=117; 15'd24815: duty=124;
15'd24816: duty=110; 15'd24817: duty=104; 15'd24818: duty=119; 15'd24819: duty=118; 15'd24820: duty=120; 15'd24821: duty=127; 15'd24822: duty=140; 15'd24823: duty=145;
15'd24824: duty=132; 15'd24825: duty=136; 15'd24826: duty=145; 15'd24827: duty=144; 15'd24828: duty=140; 15'd24829: duty=142; 15'd24830: duty=131; 15'd24831: duty=136;
15'd24832: duty=143; 15'd24833: duty=142; 15'd24834: duty=157; 15'd24835: duty=165; 15'd24836: duty=153; 15'd24837: duty=157; 15'd24838: duty=170; 15'd24839: duty=165;
15'd24840: duty=169; 15'd24841: duty=164; 15'd24842: duty=157; 15'd24843: duty=158; 15'd24844: duty=158; 15'd24845: duty=158; 15'd24846: duty=162; 15'd24847: duty=161;
15'd24848: duty=155; 15'd24849: duty=148; 15'd24850: duty=152; 15'd24851: duty=150; 15'd24852: duty=155; 15'd24853: duty=159; 15'd24854: duty=143; 15'd24855: duty=137;
15'd24856: duty=139; 15'd24857: duty=146; 15'd24858: duty=137; 15'd24859: duty=131; 15'd24860: duty=133; 15'd24861: duty=123; 15'd24862: duty=133; 15'd24863: duty=130;
15'd24864: duty=118; 15'd24865: duty=115; 15'd24866: duty=109; 15'd24867: duty=124; 15'd24868: duty=115; 15'd24869: duty=110; 15'd24870: duty=120; 15'd24871: duty=105;
15'd24872: duty=108; 15'd24873: duty=98; 15'd24874: duty=93; 15'd24875: duty=115; 15'd24876: duty=102; 15'd24877: duty=111; 15'd24878: duty=104; 15'd24879: duty=101;
15'd24880: duty=104; 15'd24881: duty=105; 15'd24882: duty=104; 15'd24883: duty=105; 15'd24884: duty=107; 15'd24885: duty=110; 15'd24886: duty=120; 15'd24887: duty=115;
15'd24888: duty=120; 15'd24889: duty=124; 15'd24890: duty=119; 15'd24891: duty=117; 15'd24892: duty=125; 15'd24893: duty=127; 15'd24894: duty=127; 15'd24895: duty=125;
15'd24896: duty=127; 15'd24897: duty=134; 15'd24898: duty=131; 15'd24899: duty=125; 15'd24900: duty=140; 15'd24901: duty=145; 15'd24902: duty=141; 15'd24903: duty=140;
15'd24904: duty=150; 15'd24905: duty=148; 15'd24906: duty=145; 15'd24907: duty=148; 15'd24908: duty=148; 15'd24909: duty=145; 15'd24910: duty=143; 15'd24911: duty=137;
15'd24912: duty=140; 15'd24913: duty=150; 15'd24914: duty=151; 15'd24915: duty=150; 15'd24916: duty=149; 15'd24917: duty=154; 15'd24918: duty=153; 15'd24919: duty=151;
15'd24920: duty=153; 15'd24921: duty=158; 15'd24922: duty=139; 15'd24923: duty=143; 15'd24924: duty=141; 15'd24925: duty=135; 15'd24926: duty=134; 15'd24927: duty=134;
15'd24928: duty=139; 15'd24929: duty=137; 15'd24930: duty=139; 15'd24931: duty=136; 15'd24932: duty=132; 15'd24933: duty=141; 15'd24934: duty=140; 15'd24935: duty=137;
15'd24936: duty=124; 15'd24937: duty=126; 15'd24938: duty=122; 15'd24939: duty=121; 15'd24940: duty=127; 15'd24941: duty=118; 15'd24942: duty=124; 15'd24943: duty=116;
15'd24944: duty=105; 15'd24945: duty=115; 15'd24946: duty=115; 15'd24947: duty=110; 15'd24948: duty=111; 15'd24949: duty=108; 15'd24950: duty=107; 15'd24951: duty=113;
15'd24952: duty=124; 15'd24953: duty=118; 15'd24954: duty=116; 15'd24955: duty=108; 15'd24956: duty=119; 15'd24957: duty=124; 15'd24958: duty=113; 15'd24959: duty=116;
15'd24960: duty=124; 15'd24961: duty=119; 15'd24962: duty=124; 15'd24963: duty=129; 15'd24964: duty=123; 15'd24965: duty=122; 15'd24966: duty=123; 15'd24967: duty=125;
15'd24968: duty=130; 15'd24969: duty=127; 15'd24970: duty=128; 15'd24971: duty=132; 15'd24972: duty=135; 15'd24973: duty=140; 15'd24974: duty=136; 15'd24975: duty=141;
15'd24976: duty=144; 15'd24977: duty=148; 15'd24978: duty=142; 15'd24979: duty=144; 15'd24980: duty=146; 15'd24981: duty=140; 15'd24982: duty=131; 15'd24983: duty=140;
15'd24984: duty=141; 15'd24985: duty=138; 15'd24986: duty=147; 15'd24987: duty=151; 15'd24988: duty=152; 15'd24989: duty=151; 15'd24990: duty=148; 15'd24991: duty=146;
15'd24992: duty=144; 15'd24993: duty=143; 15'd24994: duty=145; 15'd24995: duty=142; 15'd24996: duty=139; 15'd24997: duty=134; 15'd24998: duty=131; 15'd24999: duty=131;
15'd25000: duty=137; 15'd25001: duty=140; 15'd25002: duty=139; 15'd25003: duty=136; 15'd25004: duty=136; 15'd25005: duty=141; 15'd25006: duty=142; 15'd25007: duty=137;
15'd25008: duty=134; 15'd25009: duty=130; 15'd25010: duty=124; 15'd25011: duty=124; 15'd25012: duty=118; 15'd25013: duty=123; 15'd25014: duty=116; 15'd25015: duty=110;
15'd25016: duty=116; 15'd25017: duty=112; 15'd25018: duty=119; 15'd25019: duty=121; 15'd25020: duty=113; 15'd25021: duty=104; 15'd25022: duty=108; 15'd25023: duty=105;
15'd25024: duty=110; 15'd25025: duty=115; 15'd25026: duty=108; 15'd25027: duty=121; 15'd25028: duty=116; 15'd25029: duty=118; 15'd25030: duty=129; 15'd25031: duty=125;
15'd25032: duty=124; 15'd25033: duty=124; 15'd25034: duty=129; 15'd25035: duty=121; 15'd25036: duty=118; 15'd25037: duty=118; 15'd25038: duty=121; 15'd25039: duty=124;
15'd25040: duty=130; 15'd25041: duty=141; 15'd25042: duty=145; 15'd25043: duty=142; 15'd25044: duty=136; 15'd25045: duty=128; 15'd25046: duty=132; 15'd25047: duty=143;
15'd25048: duty=140; 15'd25049: duty=134; 15'd25050: duty=140; 15'd25051: duty=145; 15'd25052: duty=148; 15'd25053: duty=145; 15'd25054: duty=149; 15'd25055: duty=149;
15'd25056: duty=138; 15'd25057: duty=136; 15'd25058: duty=140; 15'd25059: duty=140; 15'd25060: duty=134; 15'd25061: duty=137; 15'd25062: duty=139; 15'd25063: duty=142;
15'd25064: duty=146; 15'd25065: duty=151; 15'd25066: duty=153; 15'd25067: duty=151; 15'd25068: duty=140; 15'd25069: duty=148; 15'd25070: duty=151; 15'd25071: duty=143;
15'd25072: duty=137; 15'd25073: duty=137; 15'd25074: duty=139; 15'd25075: duty=136; 15'd25076: duty=138; 15'd25077: duty=142; 15'd25078: duty=134; 15'd25079: duty=127;
15'd25080: duty=131; 15'd25081: duty=128; 15'd25082: duty=126; 15'd25083: duty=131; 15'd25084: duty=119; 15'd25085: duty=114; 15'd25086: duty=115; 15'd25087: duty=98;
15'd25088: duty=107; 15'd25089: duty=118; 15'd25090: duty=121; 15'd25091: duty=114; 15'd25092: duty=121; 15'd25093: duty=116; 15'd25094: duty=116; 15'd25095: duty=116;
15'd25096: duty=126; 15'd25097: duty=110; 15'd25098: duty=107; 15'd25099: duty=115; 15'd25100: duty=116; 15'd25101: duty=122; 15'd25102: duty=104; 15'd25103: duty=102;
15'd25104: duty=104; 15'd25105: duty=111; 15'd25106: duty=119; 15'd25107: duty=122; 15'd25108: duty=122; 15'd25109: duty=127; 15'd25110: duty=131; 15'd25111: duty=129;
15'd25112: duty=119; 15'd25113: duty=127; 15'd25114: duty=131; 15'd25115: duty=128; 15'd25116: duty=130; 15'd25117: duty=134; 15'd25118: duty=134; 15'd25119: duty=128;
15'd25120: duty=122; 15'd25121: duty=133; 15'd25122: duty=136; 15'd25123: duty=139; 15'd25124: duty=142; 15'd25125: duty=140; 15'd25126: duty=146; 15'd25127: duty=148;
15'd25128: duty=145; 15'd25129: duty=151; 15'd25130: duty=144; 15'd25131: duty=131; 15'd25132: duty=142; 15'd25133: duty=142; 15'd25134: duty=153; 15'd25135: duty=154;
15'd25136: duty=153; 15'd25137: duty=159; 15'd25138: duty=156; 15'd25139: duty=154; 15'd25140: duty=160; 15'd25141: duty=166; 15'd25142: duty=164; 15'd25143: duty=163;
15'd25144: duty=159; 15'd25145: duty=156; 15'd25146: duty=148; 15'd25147: duty=148; 15'd25148: duty=144; 15'd25149: duty=136; 15'd25150: duty=139; 15'd25151: duty=143;
15'd25152: duty=138; 15'd25153: duty=137; 15'd25154: duty=134; 15'd25155: duty=132; 15'd25156: duty=130; 15'd25157: duty=111; 15'd25158: duty=128; 15'd25159: duty=125;
15'd25160: duty=123; 15'd25161: duty=117; 15'd25162: duty=118; 15'd25163: duty=116; 15'd25164: duty=109; 15'd25165: duty=109; 15'd25166: duty=103; 15'd25167: duty=113;
15'd25168: duty=104; 15'd25169: duty=116; 15'd25170: duty=104; 15'd25171: duty=99; 15'd25172: duty=100; 15'd25173: duty=87; 15'd25174: duty=94; 15'd25175: duty=96;
15'd25176: duty=101; 15'd25177: duty=100; 15'd25178: duty=101; 15'd25179: duty=107; 15'd25180: duty=120; 15'd25181: duty=118; 15'd25182: duty=121; 15'd25183: duty=129;
15'd25184: duty=118; 15'd25185: duty=125; 15'd25186: duty=123; 15'd25187: duty=119; 15'd25188: duty=103; 15'd25189: duty=105; 15'd25190: duty=111; 15'd25191: duty=118;
15'd25192: duty=133; 15'd25193: duty=128; 15'd25194: duty=127; 15'd25195: duty=134; 15'd25196: duty=137; 15'd25197: duty=142; 15'd25198: duty=142; 15'd25199: duty=149;
15'd25200: duty=148; 15'd25201: duty=139; 15'd25202: duty=139; 15'd25203: duty=142; 15'd25204: duty=153; 15'd25205: duty=148; 15'd25206: duty=150; 15'd25207: duty=146;
15'd25208: duty=156; 15'd25209: duty=156; 15'd25210: duty=148; 15'd25211: duty=151; 15'd25212: duty=146; 15'd25213: duty=159; 15'd25214: duty=162; 15'd25215: duty=163;
15'd25216: duty=165; 15'd25217: duty=165; 15'd25218: duty=168; 15'd25219: duty=165; 15'd25220: duty=162; 15'd25221: duty=153; 15'd25222: duty=153; 15'd25223: duty=150;
15'd25224: duty=149; 15'd25225: duty=143; 15'd25226: duty=139; 15'd25227: duty=145; 15'd25228: duty=136; 15'd25229: duty=136; 15'd25230: duty=130; 15'd25231: duty=136;
15'd25232: duty=134; 15'd25233: duty=134; 15'd25234: duty=125; 15'd25235: duty=119; 15'd25236: duty=122; 15'd25237: duty=112; 15'd25238: duty=121; 15'd25239: duty=116;
15'd25240: duty=119; 15'd25241: duty=113; 15'd25242: duty=110; 15'd25243: duty=118; 15'd25244: duty=119; 15'd25245: duty=96; 15'd25246: duty=99; 15'd25247: duty=109;
15'd25248: duty=105; 15'd25249: duty=113; 15'd25250: duty=100; 15'd25251: duty=111; 15'd25252: duty=104; 15'd25253: duty=102; 15'd25254: duty=105; 15'd25255: duty=116;
15'd25256: duty=108; 15'd25257: duty=102; 15'd25258: duty=115; 15'd25259: duty=109; 15'd25260: duty=118; 15'd25261: duty=114; 15'd25262: duty=121; 15'd25263: duty=118;
15'd25264: duty=124; 15'd25265: duty=129; 15'd25266: duty=136; 15'd25267: duty=133; 15'd25268: duty=121; 15'd25269: duty=127; 15'd25270: duty=121; 15'd25271: duty=119;
15'd25272: duty=127; 15'd25273: duty=134; 15'd25274: duty=137; 15'd25275: duty=143; 15'd25276: duty=153; 15'd25277: duty=165; 15'd25278: duty=161; 15'd25279: duty=153;
15'd25280: duty=144; 15'd25281: duty=145; 15'd25282: duty=142; 15'd25283: duty=149; 15'd25284: duty=151; 15'd25285: duty=152; 15'd25286: duty=154; 15'd25287: duty=143;
15'd25288: duty=151; 15'd25289: duty=154; 15'd25290: duty=156; 15'd25291: duty=157; 15'd25292: duty=159; 15'd25293: duty=148; 15'd25294: duty=142; 15'd25295: duty=149;
15'd25296: duty=143; 15'd25297: duty=142; 15'd25298: duty=141; 15'd25299: duty=152; 15'd25300: duty=153; 15'd25301: duty=143; 15'd25302: duty=140; 15'd25303: duty=151;
15'd25304: duty=140; 15'd25305: duty=129; 15'd25306: duty=139; 15'd25307: duty=125; 15'd25308: duty=127; 15'd25309: duty=117; 15'd25310: duty=122; 15'd25311: duty=127;
15'd25312: duty=109; 15'd25313: duty=108; 15'd25314: duty=116; 15'd25315: duty=116; 15'd25316: duty=111; 15'd25317: duty=112; 15'd25318: duty=112; 15'd25319: duty=114;
15'd25320: duty=101; 15'd25321: duty=108; 15'd25322: duty=110; 15'd25323: duty=105; 15'd25324: duty=108; 15'd25325: duty=113; 15'd25326: duty=119; 15'd25327: duty=113;
15'd25328: duty=106; 15'd25329: duty=115; 15'd25330: duty=113; 15'd25331: duty=110; 15'd25332: duty=114; 15'd25333: duty=113; 15'd25334: duty=116; 15'd25335: duty=122;
15'd25336: duty=118; 15'd25337: duty=116; 15'd25338: duty=127; 15'd25339: duty=119; 15'd25340: duty=127; 15'd25341: duty=134; 15'd25342: duty=128; 15'd25343: duty=134;
15'd25344: duty=131; 15'd25345: duty=128; 15'd25346: duty=131; 15'd25347: duty=131; 15'd25348: duty=137; 15'd25349: duty=137; 15'd25350: duty=136; 15'd25351: duty=142;
15'd25352: duty=156; 15'd25353: duty=157; 15'd25354: duty=153; 15'd25355: duty=149; 15'd25356: duty=144; 15'd25357: duty=147; 15'd25358: duty=158; 15'd25359: duty=153;
15'd25360: duty=150; 15'd25361: duty=140; 15'd25362: duty=137; 15'd25363: duty=140; 15'd25364: duty=141; 15'd25365: duty=149; 15'd25366: duty=143; 15'd25367: duty=154;
15'd25368: duty=156; 15'd25369: duty=151; 15'd25370: duty=153; 15'd25371: duty=152; 15'd25372: duty=142; 15'd25373: duty=139; 15'd25374: duty=144; 15'd25375: duty=136;
15'd25376: duty=134; 15'd25377: duty=142; 15'd25378: duty=138; 15'd25379: duty=132; 15'd25380: duty=131; 15'd25381: duty=128; 15'd25382: duty=128; 15'd25383: duty=125;
15'd25384: duty=127; 15'd25385: duty=128; 15'd25386: duty=124; 15'd25387: duty=128; 15'd25388: duty=121; 15'd25389: duty=121; 15'd25390: duty=125; 15'd25391: duty=126;
15'd25392: duty=110; 15'd25393: duty=116; 15'd25394: duty=107; 15'd25395: duty=102; 15'd25396: duty=115; 15'd25397: duty=107; 15'd25398: duty=125; 15'd25399: duty=116;
15'd25400: duty=114; 15'd25401: duty=106; 15'd25402: duty=101; 15'd25403: duty=106; 15'd25404: duty=108; 15'd25405: duty=117; 15'd25406: duty=104; 15'd25407: duty=101;
15'd25408: duty=99; 15'd25409: duty=103; 15'd25410: duty=116; 15'd25411: duty=121; 15'd25412: duty=123; 15'd25413: duty=109; 15'd25414: duty=117; 15'd25415: duty=124;
15'd25416: duty=120; 15'd25417: duty=126; 15'd25418: duty=125; 15'd25419: duty=118; 15'd25420: duty=121; 15'd25421: duty=128; 15'd25422: duty=137; 15'd25423: duty=138;
15'd25424: duty=137; 15'd25425: duty=153; 15'd25426: duty=146; 15'd25427: duty=151; 15'd25428: duty=159; 15'd25429: duty=156; 15'd25430: duty=148; 15'd25431: duty=145;
15'd25432: duty=145; 15'd25433: duty=150; 15'd25434: duty=148; 15'd25435: duty=141; 15'd25436: duty=150; 15'd25437: duty=154; 15'd25438: duty=153; 15'd25439: duty=165;
15'd25440: duty=168; 15'd25441: duty=165; 15'd25442: duty=171; 15'd25443: duty=170; 15'd25444: duty=168; 15'd25445: duty=167; 15'd25446: duty=154; 15'd25447: duty=149;
15'd25448: duty=157; 15'd25449: duty=148; 15'd25450: duty=148; 15'd25451: duty=145; 15'd25452: duty=134; 15'd25453: duty=139; 15'd25454: duty=133; 15'd25455: duty=129;
15'd25456: duty=139; 15'd25457: duty=137; 15'd25458: duty=137; 15'd25459: duty=134; 15'd25460: duty=117; 15'd25461: duty=116; 15'd25462: duty=120; 15'd25463: duty=107;
15'd25464: duty=117; 15'd25465: duty=111; 15'd25466: duty=101; 15'd25467: duty=119; 15'd25468: duty=128; 15'd25469: duty=117; 15'd25470: duty=115; 15'd25471: duty=101;
15'd25472: duty=83; 15'd25473: duty=96; 15'd25474: duty=96; 15'd25475: duty=111; 15'd25476: duty=98; 15'd25477: duty=87; 15'd25478: duty=98; 15'd25479: duty=101;
15'd25480: duty=97; 15'd25481: duty=103; 15'd25482: duty=104; 15'd25483: duty=97; 15'd25484: duty=98; 15'd25485: duty=109; 15'd25486: duty=121; 15'd25487: duty=126;
15'd25488: duty=124; 15'd25489: duty=116; 15'd25490: duty=120; 15'd25491: duty=117; 15'd25492: duty=120; 15'd25493: duty=127; 15'd25494: duty=125; 15'd25495: duty=125;
15'd25496: duty=128; 15'd25497: duty=137; 15'd25498: duty=144; 15'd25499: duty=143; 15'd25500: duty=138; 15'd25501: duty=137; 15'd25502: duty=148; 15'd25503: duty=161;
15'd25504: duty=167; 15'd25505: duty=160; 15'd25506: duty=158; 15'd25507: duty=152; 15'd25508: duty=155; 15'd25509: duty=146; 15'd25510: duty=155; 15'd25511: duty=161;
15'd25512: duty=148; 15'd25513: duty=156; 15'd25514: duty=164; 15'd25515: duty=171; 15'd25516: duty=168; 15'd25517: duty=169; 15'd25518: duty=168; 15'd25519: duty=165;
15'd25520: duty=158; 15'd25521: duty=153; 15'd25522: duty=144; 15'd25523: duty=135; 15'd25524: duty=133; 15'd25525: duty=137; 15'd25526: duty=139; 15'd25527: duty=140;
15'd25528: duty=138; 15'd25529: duty=142; 15'd25530: duty=136; 15'd25531: duty=143; 15'd25532: duty=133; 15'd25533: duty=139; 15'd25534: duty=134; 15'd25535: duty=122;
15'd25536: duty=127; 15'd25537: duty=127; 15'd25538: duty=128; 15'd25539: duty=108; 15'd25540: duty=121; 15'd25541: duty=107; 15'd25542: duty=107; 15'd25543: duty=102;
15'd25544: duty=102; 15'd25545: duty=108; 15'd25546: duty=101; 15'd25547: duty=104; 15'd25548: duty=101; 15'd25549: duty=107; 15'd25550: duty=110; 15'd25551: duty=105;
15'd25552: duty=98; 15'd25553: duty=101; 15'd25554: duty=98; 15'd25555: duty=91; 15'd25556: duty=100; 15'd25557: duty=104; 15'd25558: duty=109; 15'd25559: duty=115;
15'd25560: duty=113; 15'd25561: duty=124; 15'd25562: duty=122; 15'd25563: duty=124; 15'd25564: duty=127; 15'd25565: duty=116; 15'd25566: duty=121; 15'd25567: duty=114;
15'd25568: duty=101; 15'd25569: duty=113; 15'd25570: duty=115; 15'd25571: duty=125; 15'd25572: duty=131; 15'd25573: duty=136; 15'd25574: duty=134; 15'd25575: duty=144;
15'd25576: duty=148; 15'd25577: duty=153; 15'd25578: duty=160; 15'd25579: duty=144; 15'd25580: duty=150; 15'd25581: duty=145; 15'd25582: duty=148; 15'd25583: duty=146;
15'd25584: duty=154; 15'd25585: duty=154; 15'd25586: duty=157; 15'd25587: duty=162; 15'd25588: duty=157; 15'd25589: duty=163; 15'd25590: duty=159; 15'd25591: duty=163;
15'd25592: duty=157; 15'd25593: duty=162; 15'd25594: duty=165; 15'd25595: duty=160; 15'd25596: duty=154; 15'd25597: duty=151; 15'd25598: duty=157; 15'd25599: duty=148;
15'd25600: duty=145; 15'd25601: duty=145; 15'd25602: duty=147; 15'd25603: duty=147; 15'd25604: duty=144; 15'd25605: duty=139; 15'd25606: duty=141; 15'd25607: duty=133;
15'd25608: duty=123; 15'd25609: duty=129; 15'd25610: duty=118; 15'd25611: duty=119; 15'd25612: duty=120; 15'd25613: duty=119; 15'd25614: duty=115; 15'd25615: duty=108;
15'd25616: duty=113; 15'd25617: duty=104; 15'd25618: duty=101; 15'd25619: duty=108; 15'd25620: duty=115; 15'd25621: duty=113; 15'd25622: duty=115; 15'd25623: duty=116;
15'd25624: duty=103; 15'd25625: duty=100; 15'd25626: duty=102; 15'd25627: duty=96; 15'd25628: duty=98; 15'd25629: duty=95; 15'd25630: duty=98; 15'd25631: duty=105;
15'd25632: duty=102; 15'd25633: duty=108; 15'd25634: duty=104; 15'd25635: duty=96; 15'd25636: duty=96; 15'd25637: duty=110; 15'd25638: duty=116; 15'd25639: duty=118;
15'd25640: duty=128; 15'd25641: duty=125; 15'd25642: duty=126; 15'd25643: duty=128; 15'd25644: duty=131; 15'd25645: duty=136; 15'd25646: duty=131; 15'd25647: duty=142;
15'd25648: duty=157; 15'd25649: duty=154; 15'd25650: duty=150; 15'd25651: duty=148; 15'd25652: duty=151; 15'd25653: duty=153; 15'd25654: duty=154; 15'd25655: duty=146;
15'd25656: duty=139; 15'd25657: duty=142; 15'd25658: duty=141; 15'd25659: duty=152; 15'd25660: duty=150; 15'd25661: duty=149; 15'd25662: duty=156; 15'd25663: duty=157;
15'd25664: duty=161; 15'd25665: duty=160; 15'd25666: duty=158; 15'd25667: duty=155; 15'd25668: duty=152; 15'd25669: duty=143; 15'd25670: duty=153; 15'd25671: duty=165;
15'd25672: duty=164; 15'd25673: duty=158; 15'd25674: duty=152; 15'd25675: duty=155; 15'd25676: duty=150; 15'd25677: duty=149; 15'd25678: duty=141; 15'd25679: duty=140;
15'd25680: duty=133; 15'd25681: duty=132; 15'd25682: duty=128; 15'd25683: duty=123; 15'd25684: duty=130; 15'd25685: duty=127; 15'd25686: duty=121; 15'd25687: duty=124;
15'd25688: duty=114; 15'd25689: duty=117; 15'd25690: duty=128; 15'd25691: duty=105; 15'd25692: duty=111; 15'd25693: duty=111; 15'd25694: duty=103; 15'd25695: duty=107;
15'd25696: duty=101; 15'd25697: duty=108; 15'd25698: duty=111; 15'd25699: duty=101; 15'd25700: duty=106; 15'd25701: duty=107; 15'd25702: duty=102; 15'd25703: duty=105;
15'd25704: duty=112; 15'd25705: duty=111; 15'd25706: duty=115; 15'd25707: duty=108; 15'd25708: duty=101; 15'd25709: duty=105; 15'd25710: duty=99; 15'd25711: duty=113;
15'd25712: duty=110; 15'd25713: duty=115; 15'd25714: duty=112; 15'd25715: duty=107; 15'd25716: duty=109; 15'd25717: duty=113; 15'd25718: duty=118; 15'd25719: duty=124;
15'd25720: duty=134; 15'd25721: duty=134; 15'd25722: duty=136; 15'd25723: duty=137; 15'd25724: duty=143; 15'd25725: duty=142; 15'd25726: duty=151; 15'd25727: duty=148;
15'd25728: duty=148; 15'd25729: duty=144; 15'd25730: duty=148; 15'd25731: duty=147; 15'd25732: duty=148; 15'd25733: duty=144; 15'd25734: duty=137; 15'd25735: duty=154;
15'd25736: duty=158; 15'd25737: duty=167; 15'd25738: duty=170; 15'd25739: duty=177; 15'd25740: duty=167; 15'd25741: duty=163; 15'd25742: duty=166; 15'd25743: duty=162;
15'd25744: duty=159; 15'd25745: duty=161; 15'd25746: duty=160; 15'd25747: duty=154; 15'd25748: duty=153; 15'd25749: duty=146; 15'd25750: duty=156; 15'd25751: duty=154;
15'd25752: duty=139; 15'd25753: duty=149; 15'd25754: duty=137; 15'd25755: duty=137; 15'd25756: duty=137; 15'd25757: duty=134; 15'd25758: duty=136; 15'd25759: duty=122;
15'd25760: duty=122; 15'd25761: duty=125; 15'd25762: duty=124; 15'd25763: duty=115; 15'd25764: duty=119; 15'd25765: duty=115; 15'd25766: duty=115; 15'd25767: duty=120;
15'd25768: duty=110; 15'd25769: duty=96; 15'd25770: duty=98; 15'd25771: duty=90; 15'd25772: duty=98; 15'd25773: duty=102; 15'd25774: duty=115; 15'd25775: duty=115;
15'd25776: duty=100; 15'd25777: duty=105; 15'd25778: duty=96; 15'd25779: duty=108; 15'd25780: duty=99; 15'd25781: duty=108; 15'd25782: duty=106; 15'd25783: duty=110;
15'd25784: duty=118; 15'd25785: duty=110; 15'd25786: duty=113; 15'd25787: duty=113; 15'd25788: duty=118; 15'd25789: duty=111; 15'd25790: duty=118; 15'd25791: duty=121;
15'd25792: duty=124; 15'd25793: duty=121; 15'd25794: duty=124; 15'd25795: duty=127; 15'd25796: duty=118; 15'd25797: duty=125; 15'd25798: duty=126; 15'd25799: duty=140;
15'd25800: duty=136; 15'd25801: duty=139; 15'd25802: duty=150; 15'd25803: duty=139; 15'd25804: duty=139; 15'd25805: duty=136; 15'd25806: duty=142; 15'd25807: duty=139;
15'd25808: duty=136; 15'd25809: duty=136; 15'd25810: duty=140; 15'd25811: duty=148; 15'd25812: duty=156; 15'd25813: duty=165; 15'd25814: duty=162; 15'd25815: duty=162;
15'd25816: duty=157; 15'd25817: duty=159; 15'd25818: duty=168; 15'd25819: duty=165; 15'd25820: duty=160; 15'd25821: duty=150; 15'd25822: duty=149; 15'd25823: duty=152;
15'd25824: duty=148; 15'd25825: duty=145; 15'd25826: duty=137; 15'd25827: duty=133; 15'd25828: duty=137; 15'd25829: duty=140; 15'd25830: duty=147; 15'd25831: duty=148;
15'd25832: duty=150; 15'd25833: duty=145; 15'd25834: duty=136; 15'd25835: duty=137; 15'd25836: duty=132; 15'd25837: duty=133; 15'd25838: duty=134; 15'd25839: duty=125;
15'd25840: duty=131; 15'd25841: duty=128; 15'd25842: duty=119; 15'd25843: duty=121; 15'd25844: duty=116; 15'd25845: duty=110; 15'd25846: duty=107; 15'd25847: duty=105;
15'd25848: duty=93; 15'd25849: duty=93; 15'd25850: duty=104; 15'd25851: duty=104; 15'd25852: duty=105; 15'd25853: duty=99; 15'd25854: duty=101; 15'd25855: duty=109;
15'd25856: duty=109; 15'd25857: duty=112; 15'd25858: duty=128; 15'd25859: duty=131; 15'd25860: duty=117; 15'd25861: duty=115; 15'd25862: duty=113; 15'd25863: duty=112;
15'd25864: duty=112; 15'd25865: duty=118; 15'd25866: duty=115; 15'd25867: duty=114; 15'd25868: duty=110; 15'd25869: duty=112; 15'd25870: duty=115; 15'd25871: duty=116;
15'd25872: duty=128; 15'd25873: duty=131; 15'd25874: duty=137; 15'd25875: duty=136; 15'd25876: duty=136; 15'd25877: duty=139; 15'd25878: duty=131; 15'd25879: duty=137;
15'd25880: duty=142; 15'd25881: duty=133; 15'd25882: duty=128; 15'd25883: duty=145; 15'd25884: duty=134; 15'd25885: duty=139; 15'd25886: duty=149; 15'd25887: duty=154;
15'd25888: duty=154; 15'd25889: duty=148; 15'd25890: duty=152; 15'd25891: duty=150; 15'd25892: duty=160; 15'd25893: duty=158; 15'd25894: duty=165; 15'd25895: duty=153;
15'd25896: duty=156; 15'd25897: duty=155; 15'd25898: duty=152; 15'd25899: duty=145; 15'd25900: duty=146; 15'd25901: duty=139; 15'd25902: duty=143; 15'd25903: duty=142;
15'd25904: duty=146; 15'd25905: duty=145; 15'd25906: duty=139; 15'd25907: duty=144; 15'd25908: duty=129; 15'd25909: duty=135; 15'd25910: duty=125; 15'd25911: duty=135;
15'd25912: duty=119; 15'd25913: duty=118; 15'd25914: duty=137; 15'd25915: duty=123; 15'd25916: duty=111; 15'd25917: duty=121; 15'd25918: duty=107; 15'd25919: duty=109;
15'd25920: duty=110; 15'd25921: duty=112; 15'd25922: duty=122; 15'd25923: duty=119; 15'd25924: duty=116; 15'd25925: duty=113; 15'd25926: duty=113; 15'd25927: duty=106;
15'd25928: duty=113; 15'd25929: duty=113; 15'd25930: duty=125; 15'd25931: duty=128; 15'd25932: duty=119; 15'd25933: duty=115; 15'd25934: duty=121; 15'd25935: duty=107;
15'd25936: duty=105; 15'd25937: duty=115; 15'd25938: duty=119; 15'd25939: duty=126; 15'd25940: duty=121; 15'd25941: duty=123; 15'd25942: duty=119; 15'd25943: duty=126;
15'd25944: duty=128; 15'd25945: duty=125; 15'd25946: duty=139; 15'd25947: duty=128; 15'd25948: duty=136; 15'd25949: duty=136; 15'd25950: duty=131; 15'd25951: duty=140;
15'd25952: duty=137; 15'd25953: duty=132; 15'd25954: duty=133; 15'd25955: duty=140; 15'd25956: duty=138; 15'd25957: duty=148; 15'd25958: duty=149; 15'd25959: duty=154;
15'd25960: duty=156; 15'd25961: duty=152; 15'd25962: duty=156; 15'd25963: duty=155; 15'd25964: duty=153; 15'd25965: duty=157; 15'd25966: duty=156; 15'd25967: duty=153;
15'd25968: duty=150; 15'd25969: duty=144; 15'd25970: duty=136; 15'd25971: duty=135; 15'd25972: duty=132; 15'd25973: duty=141; 15'd25974: duty=147; 15'd25975: duty=146;
15'd25976: duty=152; 15'd25977: duty=150; 15'd25978: duty=150; 15'd25979: duty=147; 15'd25980: duty=143; 15'd25981: duty=144; 15'd25982: duty=144; 15'd25983: duty=132;
15'd25984: duty=127; 15'd25985: duty=126; 15'd25986: duty=116; 15'd25987: duty=117; 15'd25988: duty=135; 15'd25989: duty=128; 15'd25990: duty=116; 15'd25991: duty=126;
15'd25992: duty=112; 15'd25993: duty=114; 15'd25994: duty=123; 15'd25995: duty=119; 15'd25996: duty=125; 15'd25997: duty=117; 15'd25998: duty=126; 15'd25999: duty=123;
15'd26000: duty=123; 15'd26001: duty=105; 15'd26002: duty=106; 15'd26003: duty=105; 15'd26004: duty=91; 15'd26005: duty=104; 15'd26006: duty=98; 15'd26007: duty=114;
15'd26008: duty=113; 15'd26009: duty=111; 15'd26010: duty=112; 15'd26011: duty=116; 15'd26012: duty=118; 15'd26013: duty=117; 15'd26014: duty=118; 15'd26015: duty=112;
15'd26016: duty=109; 15'd26017: duty=106; 15'd26018: duty=112; 15'd26019: duty=126; 15'd26020: duty=125; 15'd26021: duty=136; 15'd26022: duty=143; 15'd26023: duty=136;
15'd26024: duty=132; 15'd26025: duty=138; 15'd26026: duty=140; 15'd26027: duty=133; 15'd26028: duty=128; 15'd26029: duty=132; 15'd26030: duty=134; 15'd26031: duty=131;
15'd26032: duty=136; 15'd26033: duty=139; 15'd26034: duty=152; 15'd26035: duty=153; 15'd26036: duty=159; 15'd26037: duty=157; 15'd26038: duty=152; 15'd26039: duty=151;
15'd26040: duty=151; 15'd26041: duty=149; 15'd26042: duty=147; 15'd26043: duty=151; 15'd26044: duty=143; 15'd26045: duty=143; 15'd26046: duty=148; 15'd26047: duty=151;
15'd26048: duty=148; 15'd26049: duty=143; 15'd26050: duty=145; 15'd26051: duty=146; 15'd26052: duty=147; 15'd26053: duty=141; 15'd26054: duty=145; 15'd26055: duty=148;
15'd26056: duty=139; 15'd26057: duty=129; 15'd26058: duty=130; 15'd26059: duty=140; 15'd26060: duty=123; 15'd26061: duty=122; 15'd26062: duty=126; 15'd26063: duty=119;
15'd26064: duty=123; 15'd26065: duty=122; 15'd26066: duty=112; 15'd26067: duty=111; 15'd26068: duty=115; 15'd26069: duty=114; 15'd26070: duty=120; 15'd26071: duty=116;
15'd26072: duty=120; 15'd26073: duty=122; 15'd26074: duty=111; 15'd26075: duty=112; 15'd26076: duty=115; 15'd26077: duty=113; 15'd26078: duty=117; 15'd26079: duty=111;
15'd26080: duty=114; 15'd26081: duty=125; 15'd26082: duty=111; 15'd26083: duty=118; 15'd26084: duty=126; 15'd26085: duty=132; 15'd26086: duty=132; 15'd26087: duty=124;
15'd26088: duty=133; 15'd26089: duty=133; 15'd26090: duty=124; 15'd26091: duty=127; 15'd26092: duty=131; 15'd26093: duty=129; 15'd26094: duty=126; 15'd26095: duty=134;
15'd26096: duty=133; 15'd26097: duty=131; 15'd26098: duty=130; 15'd26099: duty=129; 15'd26100: duty=139; 15'd26101: duty=137; 15'd26102: duty=136; 15'd26103: duty=134;
15'd26104: duty=134; 15'd26105: duty=140; 15'd26106: duty=135; 15'd26107: duty=131; 15'd26108: duty=134; 15'd26109: duty=137; 15'd26110: duty=153; 15'd26111: duty=153;
15'd26112: duty=158; 15'd26113: duty=154; 15'd26114: duty=155; 15'd26115: duty=149; 15'd26116: duty=145; 15'd26117: duty=154; 15'd26118: duty=140; 15'd26119: duty=133;
15'd26120: duty=130; 15'd26121: duty=133; 15'd26122: duty=128; 15'd26123: duty=135; 15'd26124: duty=134; 15'd26125: duty=136; 15'd26126: duty=134; 15'd26127: duty=139;
15'd26128: duty=131; 15'd26129: duty=143; 15'd26130: duty=139; 15'd26131: duty=112; 15'd26132: duty=125; 15'd26133: duty=115; 15'd26134: duty=118; 15'd26135: duty=118;
15'd26136: duty=119; 15'd26137: duty=128; 15'd26138: duty=133; 15'd26139: duty=140; 15'd26140: duty=133; 15'd26141: duty=127; 15'd26142: duty=121; 15'd26143: duty=119;
15'd26144: duty=121; 15'd26145: duty=111; 15'd26146: duty=115; 15'd26147: duty=114; 15'd26148: duty=110; 15'd26149: duty=111; 15'd26150: duty=121; 15'd26151: duty=123;
15'd26152: duty=120; 15'd26153: duty=117; 15'd26154: duty=120; 15'd26155: duty=132; 15'd26156: duty=131; 15'd26157: duty=132; 15'd26158: duty=127; 15'd26159: duty=127;
15'd26160: duty=130; 15'd26161: duty=134; 15'd26162: duty=132; 15'd26163: duty=132; 15'd26164: duty=120; 15'd26165: duty=113; 15'd26166: duty=121; 15'd26167: duty=125;
15'd26168: duty=133; 15'd26169: duty=134; 15'd26170: duty=133; 15'd26171: duty=145; 15'd26172: duty=149; 15'd26173: duty=146; 15'd26174: duty=147; 15'd26175: duty=143;
15'd26176: duty=138; 15'd26177: duty=132; 15'd26178: duty=135; 15'd26179: duty=132; 15'd26180: duty=135; 15'd26181: duty=141; 15'd26182: duty=135; 15'd26183: duty=140;
15'd26184: duty=144; 15'd26185: duty=151; 15'd26186: duty=152; 15'd26187: duty=155; 15'd26188: duty=149; 15'd26189: duty=140; 15'd26190: duty=145; 15'd26191: duty=142;
15'd26192: duty=139; 15'd26193: duty=138; 15'd26194: duty=139; 15'd26195: duty=132; 15'd26196: duty=123; 15'd26197: duty=134; 15'd26198: duty=139; 15'd26199: duty=140;
15'd26200: duty=137; 15'd26201: duty=131; 15'd26202: duty=123; 15'd26203: duty=117; 15'd26204: duty=120; 15'd26205: duty=116; 15'd26206: duty=118; 15'd26207: duty=113;
15'd26208: duty=113; 15'd26209: duty=113; 15'd26210: duty=115; 15'd26211: duty=113; 15'd26212: duty=110; 15'd26213: duty=111; 15'd26214: duty=110; 15'd26215: duty=108;
15'd26216: duty=113; 15'd26217: duty=121; 15'd26218: duty=108; 15'd26219: duty=110; 15'd26220: duty=112; 15'd26221: duty=102; 15'd26222: duty=110; 15'd26223: duty=113;
15'd26224: duty=112; 15'd26225: duty=115; 15'd26226: duty=119; 15'd26227: duty=130; 15'd26228: duty=131; 15'd26229: duty=130; 15'd26230: duty=128; 15'd26231: duty=131;
15'd26232: duty=128; 15'd26233: duty=133; 15'd26234: duty=138; 15'd26235: duty=136; 15'd26236: duty=133; 15'd26237: duty=139; 15'd26238: duty=144; 15'd26239: duty=140;
15'd26240: duty=136; 15'd26241: duty=141; 15'd26242: duty=140; 15'd26243: duty=142; 15'd26244: duty=151; 15'd26245: duty=151; 15'd26246: duty=153; 15'd26247: duty=139;
15'd26248: duty=142; 15'd26249: duty=150; 15'd26250: duty=148; 15'd26251: duty=141; 15'd26252: duty=148; 15'd26253: duty=148; 15'd26254: duty=151; 15'd26255: duty=156;
15'd26256: duty=152; 15'd26257: duty=160; 15'd26258: duty=155; 15'd26259: duty=154; 15'd26260: duty=156; 15'd26261: duty=151; 15'd26262: duty=153; 15'd26263: duty=150;
15'd26264: duty=142; 15'd26265: duty=145; 15'd26266: duty=146; 15'd26267: duty=144; 15'd26268: duty=145; 15'd26269: duty=142; 15'd26270: duty=134; 15'd26271: duty=137;
15'd26272: duty=130; 15'd26273: duty=137; 15'd26274: duty=139; 15'd26275: duty=121; 15'd26276: duty=118; 15'd26277: duty=110; 15'd26278: duty=118; 15'd26279: duty=116;
15'd26280: duty=123; 15'd26281: duty=121; 15'd26282: duty=115; 15'd26283: duty=118; 15'd26284: duty=114; 15'd26285: duty=119; 15'd26286: duty=107; 15'd26287: duty=113;
15'd26288: duty=115; 15'd26289: duty=107; 15'd26290: duty=109; 15'd26291: duty=111; 15'd26292: duty=117; 15'd26293: duty=111; 15'd26294: duty=107; 15'd26295: duty=96;
15'd26296: duty=104; 15'd26297: duty=96; 15'd26298: duty=93; 15'd26299: duty=110; 15'd26300: duty=107; 15'd26301: duty=113; 15'd26302: duty=106; 15'd26303: duty=109;
15'd26304: duty=113; 15'd26305: duty=119; 15'd26306: duty=121; 15'd26307: duty=118; 15'd26308: duty=125; 15'd26309: duty=124; 15'd26310: duty=122; 15'd26311: duty=114;
15'd26312: duty=116; 15'd26313: duty=116; 15'd26314: duty=118; 15'd26315: duty=119; 15'd26316: duty=119; 15'd26317: duty=136; 15'd26318: duty=136; 15'd26319: duty=148;
15'd26320: duty=145; 15'd26321: duty=139; 15'd26322: duty=145; 15'd26323: duty=143; 15'd26324: duty=148; 15'd26325: duty=151; 15'd26326: duty=145; 15'd26327: duty=143;
15'd26328: duty=150; 15'd26329: duty=151; 15'd26330: duty=166; 15'd26331: duty=164; 15'd26332: duty=166; 15'd26333: duty=171; 15'd26334: duty=163; 15'd26335: duty=166;
15'd26336: duty=164; 15'd26337: duty=163; 15'd26338: duty=162; 15'd26339: duty=158; 15'd26340: duty=158; 15'd26341: duty=155; 15'd26342: duty=149; 15'd26343: duty=148;
15'd26344: duty=147; 15'd26345: duty=138; 15'd26346: duty=145; 15'd26347: duty=144; 15'd26348: duty=136; 15'd26349: duty=138; 15'd26350: duty=136; 15'd26351: duty=137;
15'd26352: duty=129; 15'd26353: duty=122; 15'd26354: duty=130; 15'd26355: duty=126; 15'd26356: duty=112; 15'd26357: duty=120; 15'd26358: duty=124; 15'd26359: duty=125;
15'd26360: duty=127; 15'd26361: duty=119; 15'd26362: duty=115; 15'd26363: duty=113; 15'd26364: duty=98; 15'd26365: duty=108; 15'd26366: duty=114; 15'd26367: duty=110;
15'd26368: duty=101; 15'd26369: duty=103; 15'd26370: duty=107; 15'd26371: duty=100; 15'd26372: duty=107; 15'd26373: duty=107; 15'd26374: duty=106; 15'd26375: duty=105;
15'd26376: duty=113; 15'd26377: duty=114; 15'd26378: duty=114; 15'd26379: duty=117; 15'd26380: duty=123; 15'd26381: duty=125; 15'd26382: duty=123; 15'd26383: duty=125;
15'd26384: duty=123; 15'd26385: duty=119; 15'd26386: duty=127; 15'd26387: duty=127; 15'd26388: duty=130; 15'd26389: duty=129; 15'd26390: duty=130; 15'd26391: duty=138;
15'd26392: duty=138; 15'd26393: duty=143; 15'd26394: duty=138; 15'd26395: duty=143; 15'd26396: duty=150; 15'd26397: duty=154; 15'd26398: duty=149; 15'd26399: duty=138;
15'd26400: duty=142; 15'd26401: duty=140; 15'd26402: duty=136; 15'd26403: duty=146; 15'd26404: duty=144; 15'd26405: duty=146; 15'd26406: duty=149; 15'd26407: duty=151;
15'd26408: duty=164; 15'd26409: duty=163; 15'd26410: duty=163; 15'd26411: duty=152; 15'd26412: duty=144; 15'd26413: duty=150; 15'd26414: duty=147; 15'd26415: duty=137;
15'd26416: duty=147; 15'd26417: duty=145; 15'd26418: duty=135; 15'd26419: duty=140; 15'd26420: duty=130; 15'd26421: duty=136; 15'd26422: duty=139; 15'd26423: duty=141;
15'd26424: duty=138; 15'd26425: duty=135; 15'd26426: duty=141; 15'd26427: duty=128; 15'd26428: duty=124; 15'd26429: duty=126; 15'd26430: duty=117; 15'd26431: duty=113;
15'd26432: duty=118; 15'd26433: duty=113; 15'd26434: duty=128; 15'd26435: duty=122; 15'd26436: duty=107; 15'd26437: duty=105; 15'd26438: duty=98; 15'd26439: duty=99;
15'd26440: duty=112; 15'd26441: duty=116; 15'd26442: duty=109; 15'd26443: duty=114; 15'd26444: duty=100; 15'd26445: duty=91; 15'd26446: duty=98; 15'd26447: duty=104;
15'd26448: duty=112; 15'd26449: duty=115; 15'd26450: duty=107; 15'd26451: duty=115; 15'd26452: duty=119; 15'd26453: duty=124; 15'd26454: duty=124; 15'd26455: duty=116;
15'd26456: duty=108; 15'd26457: duty=115; 15'd26458: duty=128; 15'd26459: duty=127; 15'd26460: duty=133; 15'd26461: duty=126; 15'd26462: duty=128; 15'd26463: duty=134;
15'd26464: duty=134; 15'd26465: duty=144; 15'd26466: duty=156; 15'd26467: duty=156; 15'd26468: duty=157; 15'd26469: duty=159; 15'd26470: duty=156; 15'd26471: duty=148;
15'd26472: duty=145; 15'd26473: duty=140; 15'd26474: duty=136; 15'd26475: duty=137; 15'd26476: duty=140; 15'd26477: duty=148; 15'd26478: duty=153; 15'd26479: duty=154;
15'd26480: duty=157; 15'd26481: duty=157; 15'd26482: duty=165; 15'd26483: duty=165; 15'd26484: duty=163; 15'd26485: duty=159; 15'd26486: duty=145; 15'd26487: duty=148;
15'd26488: duty=139; 15'd26489: duty=142; 15'd26490: duty=142; 15'd26491: duty=142; 15'd26492: duty=145; 15'd26493: duty=146; 15'd26494: duty=136; 15'd26495: duty=144;
15'd26496: duty=146; 15'd26497: duty=128; 15'd26498: duty=139; 15'd26499: duty=131; 15'd26500: duty=126; 15'd26501: duty=126; 15'd26502: duty=124; 15'd26503: duty=131;
15'd26504: duty=130; 15'd26505: duty=125; 15'd26506: duty=126; 15'd26507: duty=121; 15'd26508: duty=108; 15'd26509: duty=105; 15'd26510: duty=107; 15'd26511: duty=104;
15'd26512: duty=116; 15'd26513: duty=112; 15'd26514: duty=107; 15'd26515: duty=102; 15'd26516: duty=105; 15'd26517: duty=102; 15'd26518: duty=93; 15'd26519: duty=101;
15'd26520: duty=102; 15'd26521: duty=110; 15'd26522: duty=116; 15'd26523: duty=119; 15'd26524: duty=116; 15'd26525: duty=110; 15'd26526: duty=106; 15'd26527: duty=105;
15'd26528: duty=107; 15'd26529: duty=113; 15'd26530: duty=116; 15'd26531: duty=120; 15'd26532: duty=127; 15'd26533: duty=122; 15'd26534: duty=123; 15'd26535: duty=131;
15'd26536: duty=128; 15'd26537: duty=132; 15'd26538: duty=124; 15'd26539: duty=132; 15'd26540: duty=130; 15'd26541: duty=129; 15'd26542: duty=141; 15'd26543: duty=135;
15'd26544: duty=132; 15'd26545: duty=140; 15'd26546: duty=144; 15'd26547: duty=143; 15'd26548: duty=148; 15'd26549: duty=148; 15'd26550: duty=156; 15'd26551: duty=154;
15'd26552: duty=146; 15'd26553: duty=157; 15'd26554: duty=162; 15'd26555: duty=154; 15'd26556: duty=153; 15'd26557: duty=160; 15'd26558: duty=166; 15'd26559: duty=161;
15'd26560: duty=164; 15'd26561: duty=166; 15'd26562: duty=158; 15'd26563: duty=157; 15'd26564: duty=164; 15'd26565: duty=152; 15'd26566: duty=150; 15'd26567: duty=152;
15'd26568: duty=150; 15'd26569: duty=146; 15'd26570: duty=142; 15'd26571: duty=149; 15'd26572: duty=139; 15'd26573: duty=141; 15'd26574: duty=133; 15'd26575: duty=141;
15'd26576: duty=136; 15'd26577: duty=116; 15'd26578: duty=115; 15'd26579: duty=111; 15'd26580: duty=117; 15'd26581: duty=120; 15'd26582: duty=120; 15'd26583: duty=114;
15'd26584: duty=118; 15'd26585: duty=103; 15'd26586: duty=111; 15'd26587: duty=125; 15'd26588: duty=125; 15'd26589: duty=128; 15'd26590: duty=114; 15'd26591: duty=105;
15'd26592: duty=97; 15'd26593: duty=85; 15'd26594: duty=84; 15'd26595: duty=94; 15'd26596: duty=97; 15'd26597: duty=100; 15'd26598: duty=108; 15'd26599: duty=119;
15'd26600: duty=115; 15'd26601: duty=120; 15'd26602: duty=118; 15'd26603: duty=125; 15'd26604: duty=113; 15'd26605: duty=111; 15'd26606: duty=120; 15'd26607: duty=119;
15'd26608: duty=121; 15'd26609: duty=117; 15'd26610: duty=121; 15'd26611: duty=121; 15'd26612: duty=129; 15'd26613: duty=132; 15'd26614: duty=133; 15'd26615: duty=135;
15'd26616: duty=134; 15'd26617: duty=134; 15'd26618: duty=140; 15'd26619: duty=136; 15'd26620: duty=133; 15'd26621: duty=129; 15'd26622: duty=139; 15'd26623: duty=134;
15'd26624: duty=139; 15'd26625: duty=148; 15'd26626: duty=150; 15'd26627: duty=148; 15'd26628: duty=151; 15'd26629: duty=168; 15'd26630: duty=159; 15'd26631: duty=163;
15'd26632: duty=162; 15'd26633: duty=160; 15'd26634: duty=157; 15'd26635: duty=153; 15'd26636: duty=157; 15'd26637: duty=145; 15'd26638: duty=143; 15'd26639: duty=148;
15'd26640: duty=153; 15'd26641: duty=154; 15'd26642: duty=148; 15'd26643: duty=157; 15'd26644: duty=150; 15'd26645: duty=149; 15'd26646: duty=133; 15'd26647: duty=134;
15'd26648: duty=137; 15'd26649: duty=121; 15'd26650: duty=136; 15'd26651: duty=131; 15'd26652: duty=128; 15'd26653: duty=119; 15'd26654: duty=127; 15'd26655: duty=127;
15'd26656: duty=121; 15'd26657: duty=127; 15'd26658: duty=118; 15'd26659: duty=122; 15'd26660: duty=106; 15'd26661: duty=108; 15'd26662: duty=108; 15'd26663: duty=108;
15'd26664: duty=112; 15'd26665: duty=120; 15'd26666: duty=112; 15'd26667: duty=104; 15'd26668: duty=113; 15'd26669: duty=113; 15'd26670: duty=114; 15'd26671: duty=102;
15'd26672: duty=106; 15'd26673: duty=109; 15'd26674: duty=117; 15'd26675: duty=117; 15'd26676: duty=126; 15'd26677: duty=124; 15'd26678: duty=120; 15'd26679: duty=125;
15'd26680: duty=115; 15'd26681: duty=121; 15'd26682: duty=124; 15'd26683: duty=122; 15'd26684: duty=126; 15'd26685: duty=128; 15'd26686: duty=116; 15'd26687: duty=128;
15'd26688: duty=133; 15'd26689: duty=134; 15'd26690: duty=139; 15'd26691: duty=132; 15'd26692: duty=139; 15'd26693: duty=140; 15'd26694: duty=135; 15'd26695: duty=134;
15'd26696: duty=133; 15'd26697: duty=136; 15'd26698: duty=137; 15'd26699: duty=139; 15'd26700: duty=137; 15'd26701: duty=144; 15'd26702: duty=148; 15'd26703: duty=153;
15'd26704: duty=148; 15'd26705: duty=152; 15'd26706: duty=160; 15'd26707: duty=164; 15'd26708: duty=160; 15'd26709: duty=158; 15'd26710: duty=155; 15'd26711: duty=147;
15'd26712: duty=152; 15'd26713: duty=136; 15'd26714: duty=128; 15'd26715: duty=137; 15'd26716: duty=144; 15'd26717: duty=129; 15'd26718: duty=131; 15'd26719: duty=136;
15'd26720: duty=129; 15'd26721: duty=123; 15'd26722: duty=125; 15'd26723: duty=126; 15'd26724: duty=125; 15'd26725: duty=133; 15'd26726: duty=132; 15'd26727: duty=133;
15'd26728: duty=127; 15'd26729: duty=124; 15'd26730: duty=127; 15'd26731: duty=130; 15'd26732: duty=125; 15'd26733: duty=118; 15'd26734: duty=115; 15'd26735: duty=118;
15'd26736: duty=121; 15'd26737: duty=116; 15'd26738: duty=108; 15'd26739: duty=106; 15'd26740: duty=105; 15'd26741: duty=105; 15'd26742: duty=122; 15'd26743: duty=128;
15'd26744: duty=122; 15'd26745: duty=117; 15'd26746: duty=119; 15'd26747: duty=118; 15'd26748: duty=111; 15'd26749: duty=122; 15'd26750: duty=119; 15'd26751: duty=126;
15'd26752: duty=125; 15'd26753: duty=127; 15'd26754: duty=134; 15'd26755: duty=133; 15'd26756: duty=132; 15'd26757: duty=130; 15'd26758: duty=124; 15'd26759: duty=119;
15'd26760: duty=130; 15'd26761: duty=134; 15'd26762: duty=136; 15'd26763: duty=143; 15'd26764: duty=142; 15'd26765: duty=147; 15'd26766: duty=151; 15'd26767: duty=147;
15'd26768: duty=141; 15'd26769: duty=136; 15'd26770: duty=151; 15'd26771: duty=145; 15'd26772: duty=153; 15'd26773: duty=152; 15'd26774: duty=148; 15'd26775: duty=152;
15'd26776: duty=159; 15'd26777: duty=163; 15'd26778: duty=162; 15'd26779: duty=165; 15'd26780: duty=153; 15'd26781: duty=160; 15'd26782: duty=147; 15'd26783: duty=149;
15'd26784: duty=144; 15'd26785: duty=132; 15'd26786: duty=144; 15'd26787: duty=132; 15'd26788: duty=133; 15'd26789: duty=145; 15'd26790: duty=144; 15'd26791: duty=147;
15'd26792: duty=139; 15'd26793: duty=132; 15'd26794: duty=127; 15'd26795: duty=125; 15'd26796: duty=115; 15'd26797: duty=119; 15'd26798: duty=123; 15'd26799: duty=117;
15'd26800: duty=109; 15'd26801: duty=109; 15'd26802: duty=121; 15'd26803: duty=111; 15'd26804: duty=109; 15'd26805: duty=106; 15'd26806: duty=101; 15'd26807: duty=95;
15'd26808: duty=98; 15'd26809: duty=97; 15'd26810: duty=100; 15'd26811: duty=106; 15'd26812: duty=103; 15'd26813: duty=102; 15'd26814: duty=101; 15'd26815: duty=105;
15'd26816: duty=110; 15'd26817: duty=108; 15'd26818: duty=101; 15'd26819: duty=100; 15'd26820: duty=115; 15'd26821: duty=119; 15'd26822: duty=126; 15'd26823: duty=122;
15'd26824: duty=116; 15'd26825: duty=117; 15'd26826: duty=112; 15'd26827: duty=128; 15'd26828: duty=121; 15'd26829: duty=126; 15'd26830: duty=122; 15'd26831: duty=128;
15'd26832: duty=124; 15'd26833: duty=134; 15'd26834: duty=141; 15'd26835: duty=136; 15'd26836: duty=148; 15'd26837: duty=141; 15'd26838: duty=153; 15'd26839: duty=149;
15'd26840: duty=149; 15'd26841: duty=145; 15'd26842: duty=145; 15'd26843: duty=145; 15'd26844: duty=142; 15'd26845: duty=146; 15'd26846: duty=151; 15'd26847: duty=157;
15'd26848: duty=148; 15'd26849: duty=154; 15'd26850: duty=161; 15'd26851: duty=163; 15'd26852: duty=164; 15'd26853: duty=165; 15'd26854: duty=167; 15'd26855: duty=157;
15'd26856: duty=156; 15'd26857: duty=162; 15'd26858: duty=163; 15'd26859: duty=155; 15'd26860: duty=151; 15'd26861: duty=151; 15'd26862: duty=151; 15'd26863: duty=148;
15'd26864: duty=154; 15'd26865: duty=148; 15'd26866: duty=139; 15'd26867: duty=143; 15'd26868: duty=138; 15'd26869: duty=137; 15'd26870: duty=130; 15'd26871: duty=132;
15'd26872: duty=130; 15'd26873: duty=119; 15'd26874: duty=124; 15'd26875: duty=122; 15'd26876: duty=120; 15'd26877: duty=125; 15'd26878: duty=122; 15'd26879: duty=122;
15'd26880: duty=112; 15'd26881: duty=117; 15'd26882: duty=118; 15'd26883: duty=107; 15'd26884: duty=104; 15'd26885: duty=99; 15'd26886: duty=99; 15'd26887: duty=96;
15'd26888: duty=98; 15'd26889: duty=95; 15'd26890: duty=105; 15'd26891: duty=113; 15'd26892: duty=107; 15'd26893: duty=105; 15'd26894: duty=105; 15'd26895: duty=107;
15'd26896: duty=115; 15'd26897: duty=118; 15'd26898: duty=111; 15'd26899: duty=124; 15'd26900: duty=113; 15'd26901: duty=107; 15'd26902: duty=110; 15'd26903: duty=116;
15'd26904: duty=129; 15'd26905: duty=128; 15'd26906: duty=119; 15'd26907: duty=118; 15'd26908: duty=130; 15'd26909: duty=134; 15'd26910: duty=146; 15'd26911: duty=142;
15'd26912: duty=129; 15'd26913: duty=133; 15'd26914: duty=145; 15'd26915: duty=139; 15'd26916: duty=131; 15'd26917: duty=134; 15'd26918: duty=133; 15'd26919: duty=125;
15'd26920: duty=128; 15'd26921: duty=135; 15'd26922: duty=147; 15'd26923: duty=153; 15'd26924: duty=151; 15'd26925: duty=148; 15'd26926: duty=149; 15'd26927: duty=159;
15'd26928: duty=165; 15'd26929: duty=168; 15'd26930: duty=168; 15'd26931: duty=153; 15'd26932: duty=148; 15'd26933: duty=145; 15'd26934: duty=139; 15'd26935: duty=145;
15'd26936: duty=142; 15'd26937: duty=150; 15'd26938: duty=149; 15'd26939: duty=150; 15'd26940: duty=143; 15'd26941: duty=135; 15'd26942: duty=135; 15'd26943: duty=127;
15'd26944: duty=130; 15'd26945: duty=142; 15'd26946: duty=134; 15'd26947: duty=136; 15'd26948: duty=128; 15'd26949: duty=124; 15'd26950: duty=131; 15'd26951: duty=133;
15'd26952: duty=130; 15'd26953: duty=127; 15'd26954: duty=134; 15'd26955: duty=127; 15'd26956: duty=129; 15'd26957: duty=121; 15'd26958: duty=113; 15'd26959: duty=109;
15'd26960: duty=104; 15'd26961: duty=106; 15'd26962: duty=110; 15'd26963: duty=106; 15'd26964: duty=105; 15'd26965: duty=110; 15'd26966: duty=107; 15'd26967: duty=106;
15'd26968: duty=108; 15'd26969: duty=118; 15'd26970: duty=118; 15'd26971: duty=112; 15'd26972: duty=124; 15'd26973: duty=122; 15'd26974: duty=125; 15'd26975: duty=127;
15'd26976: duty=128; 15'd26977: duty=125; 15'd26978: duty=116; 15'd26979: duty=124; 15'd26980: duty=129; 15'd26981: duty=131; 15'd26982: duty=130; 15'd26983: duty=135;
15'd26984: duty=140; 15'd26985: duty=146; 15'd26986: duty=150; 15'd26987: duty=139; 15'd26988: duty=142; 15'd26989: duty=139; 15'd26990: duty=119; 15'd26991: duty=128;
15'd26992: duty=130; 15'd26993: duty=121; 15'd26994: duty=127; 15'd26995: duty=126; 15'd26996: duty=130; 15'd26997: duty=145; 15'd26998: duty=148; 15'd26999: duty=154;
15'd27000: duty=159; 15'd27001: duty=148; 15'd27002: duty=154; 15'd27003: duty=160; 15'd27004: duty=146; 15'd27005: duty=145; 15'd27006: duty=142; 15'd27007: duty=135;
15'd27008: duty=140; 15'd27009: duty=142; 15'd27010: duty=137; 15'd27011: duty=149; 15'd27012: duty=150; 15'd27013: duty=136; 15'd27014: duty=138; 15'd27015: duty=131;
15'd27016: duty=134; 15'd27017: duty=148; 15'd27018: duty=139; 15'd27019: duty=139; 15'd27020: duty=134; 15'd27021: duty=131; 15'd27022: duty=139; 15'd27023: duty=134;
15'd27024: duty=139; 15'd27025: duty=130; 15'd27026: duty=126; 15'd27027: duty=130; 15'd27028: duty=125; 15'd27029: duty=124; 15'd27030: duty=122; 15'd27031: duty=118;
15'd27032: duty=118; 15'd27033: duty=114; 15'd27034: duty=106; 15'd27035: duty=117; 15'd27036: duty=115; 15'd27037: duty=112; 15'd27038: duty=111; 15'd27039: duty=99;
15'd27040: duty=108; 15'd27041: duty=121; 15'd27042: duty=116; 15'd27043: duty=119; 15'd27044: duty=122; 15'd27045: duty=123; 15'd27046: duty=128; 15'd27047: duty=126;
15'd27048: duty=127; 15'd27049: duty=124; 15'd27050: duty=125; 15'd27051: duty=119; 15'd27052: duty=117; 15'd27053: duty=120; 15'd27054: duty=119; 15'd27055: duty=116;
15'd27056: duty=120; 15'd27057: duty=136; 15'd27058: duty=122; 15'd27059: duty=132; 15'd27060: duty=145; 15'd27061: duty=138; 15'd27062: duty=143; 15'd27063: duty=134;
15'd27064: duty=124; 15'd27065: duty=129; 15'd27066: duty=134; 15'd27067: duty=127; 15'd27068: duty=135; 15'd27069: duty=147; 15'd27070: duty=147; 15'd27071: duty=151;
15'd27072: duty=160; 15'd27073: duty=156; 15'd27074: duty=150; 15'd27075: duty=156; 15'd27076: duty=145; 15'd27077: duty=149; 15'd27078: duty=147; 15'd27079: duty=144;
15'd27080: duty=150; 15'd27081: duty=150; 15'd27082: duty=150; 15'd27083: duty=142; 15'd27084: duty=142; 15'd27085: duty=147; 15'd27086: duty=150; 15'd27087: duty=145;
15'd27088: duty=146; 15'd27089: duty=138; 15'd27090: duty=129; 15'd27091: duty=129; 15'd27092: duty=128; 15'd27093: duty=127; 15'd27094: duty=124; 15'd27095: duty=113;
15'd27096: duty=110; 15'd27097: duty=124; 15'd27098: duty=118; 15'd27099: duty=119; 15'd27100: duty=114; 15'd27101: duty=109; 15'd27102: duty=104; 15'd27103: duty=107;
15'd27104: duty=116; 15'd27105: duty=117; 15'd27106: duty=112; 15'd27107: duty=115; 15'd27108: duty=116; 15'd27109: duty=104; 15'd27110: duty=113; 15'd27111: duty=112;
15'd27112: duty=115; 15'd27113: duty=116; 15'd27114: duty=116; 15'd27115: duty=112; 15'd27116: duty=109; 15'd27117: duty=121; 15'd27118: duty=115; 15'd27119: duty=114;
15'd27120: duty=120; 15'd27121: duty=121; 15'd27122: duty=114; 15'd27123: duty=112; 15'd27124: duty=124; 15'd27125: duty=128; 15'd27126: duty=123; 15'd27127: duty=125;
15'd27128: duty=137; 15'd27129: duty=131; 15'd27130: duty=142; 15'd27131: duty=145; 15'd27132: duty=133; 15'd27133: duty=139; 15'd27134: duty=140; 15'd27135: duty=138;
15'd27136: duty=140; 15'd27137: duty=141; 15'd27138: duty=135; 15'd27139: duty=139; 15'd27140: duty=146; 15'd27141: duty=144; 15'd27142: duty=152; 15'd27143: duty=156;
15'd27144: duty=149; 15'd27145: duty=155; 15'd27146: duty=171; 15'd27147: duty=176; 15'd27148: duty=174; 15'd27149: duty=170; 15'd27150: duty=160; 15'd27151: duty=156;
15'd27152: duty=155; 15'd27153: duty=153; 15'd27154: duty=154; 15'd27155: duty=146; 15'd27156: duty=142; 15'd27157: duty=148; 15'd27158: duty=146; 15'd27159: duty=147;
15'd27160: duty=143; 15'd27161: duty=133; 15'd27162: duty=136; 15'd27163: duty=137; 15'd27164: duty=128; 15'd27165: duty=127; 15'd27166: duty=143; 15'd27167: duty=136;
15'd27168: duty=119; 15'd27169: duty=133; 15'd27170: duty=128; 15'd27171: duty=125; 15'd27172: duty=131; 15'd27173: duty=128; 15'd27174: duty=137; 15'd27175: duty=124;
15'd27176: duty=116; 15'd27177: duty=118; 15'd27178: duty=113; 15'd27179: duty=117; 15'd27180: duty=121; 15'd27181: duty=110; 15'd27182: duty=105; 15'd27183: duty=107;
15'd27184: duty=111; 15'd27185: duty=112; 15'd27186: duty=105; 15'd27187: duty=95; 15'd27188: duty=99; 15'd27189: duty=104; 15'd27190: duty=106; 15'd27191: duty=112;
15'd27192: duty=104; 15'd27193: duty=103; 15'd27194: duty=105; 15'd27195: duty=107; 15'd27196: duty=114; 15'd27197: duty=115; 15'd27198: duty=112; 15'd27199: duty=116;
15'd27200: duty=108; 15'd27201: duty=109; 15'd27202: duty=119; 15'd27203: duty=119; 15'd27204: duty=119; 15'd27205: duty=128; 15'd27206: duty=132; 15'd27207: duty=141;
15'd27208: duty=138; 15'd27209: duty=136; 15'd27210: duty=132; 15'd27211: duty=121; 15'd27212: duty=129; 15'd27213: duty=131; 15'd27214: duty=136; 15'd27215: duty=132;
15'd27216: duty=137; 15'd27217: duty=144; 15'd27218: duty=155; 15'd27219: duty=159; 15'd27220: duty=153; 15'd27221: duty=153; 15'd27222: duty=162; 15'd27223: duty=158;
15'd27224: duty=171; 15'd27225: duty=174; 15'd27226: duty=169; 15'd27227: duty=161; 15'd27228: duty=144; 15'd27229: duty=145; 15'd27230: duty=146; 15'd27231: duty=145;
15'd27232: duty=146; 15'd27233: duty=154; 15'd27234: duty=140; 15'd27235: duty=136; 15'd27236: duty=145; 15'd27237: duty=135; 15'd27238: duty=128; 15'd27239: duty=133;
15'd27240: duty=125; 15'd27241: duty=138; 15'd27242: duty=136; 15'd27243: duty=143; 15'd27244: duty=127; 15'd27245: duty=122; 15'd27246: duty=123; 15'd27247: duty=117;
15'd27248: duty=117; 15'd27249: duty=120; 15'd27250: duty=122; 15'd27251: duty=114; 15'd27252: duty=116; 15'd27253: duty=109; 15'd27254: duty=109; 15'd27255: duty=102;
15'd27256: duty=111; 15'd27257: duty=104; 15'd27258: duty=115; 15'd27259: duty=125; 15'd27260: duty=128; 15'd27261: duty=123; 15'd27262: duty=121; 15'd27263: duty=118;
15'd27264: duty=119; 15'd27265: duty=123; 15'd27266: duty=119; 15'd27267: duty=116; 15'd27268: duty=121; 15'd27269: duty=124; 15'd27270: duty=113; 15'd27271: duty=122;
15'd27272: duty=134; 15'd27273: duty=140; 15'd27274: duty=131; 15'd27275: duty=131; 15'd27276: duty=139; 15'd27277: duty=137; 15'd27278: duty=140; 15'd27279: duty=144;
15'd27280: duty=137; 15'd27281: duty=126; 15'd27282: duty=128; 15'd27283: duty=137; 15'd27284: duty=134; 15'd27285: duty=126; 15'd27286: duty=134; 15'd27287: duty=139;
15'd27288: duty=145; 15'd27289: duty=148; 15'd27290: duty=157; 15'd27291: duty=161; 15'd27292: duty=151; 15'd27293: duty=156; 15'd27294: duty=160; 15'd27295: duty=160;
15'd27296: duty=154; 15'd27297: duty=157; 15'd27298: duty=159; 15'd27299: duty=162; 15'd27300: duty=151; 15'd27301: duty=143; 15'd27302: duty=145; 15'd27303: duty=140;
15'd27304: duty=134; 15'd27305: duty=133; 15'd27306: duty=128; 15'd27307: duty=126; 15'd27308: duty=125; 15'd27309: duty=119; 15'd27310: duty=111; 15'd27311: duty=111;
15'd27312: duty=126; 15'd27313: duty=116; 15'd27314: duty=116; 15'd27315: duty=128; 15'd27316: duty=137; 15'd27317: duty=130; 15'd27318: duty=122; 15'd27319: duty=121;
15'd27320: duty=111; 15'd27321: duty=112; 15'd27322: duty=109; 15'd27323: duty=114; 15'd27324: duty=109; 15'd27325: duty=105; 15'd27326: duty=113; 15'd27327: duty=116;
15'd27328: duty=109; 15'd27329: duty=105; 15'd27330: duty=111; 15'd27331: duty=101; 15'd27332: duty=112; 15'd27333: duty=110; 15'd27334: duty=111; 15'd27335: duty=112;
15'd27336: duty=113; 15'd27337: duty=112; 15'd27338: duty=109; 15'd27339: duty=110; 15'd27340: duty=114; 15'd27341: duty=125; 15'd27342: duty=131; 15'd27343: duty=127;
15'd27344: duty=126; 15'd27345: duty=130; 15'd27346: duty=129; 15'd27347: duty=141; 15'd27348: duty=133; 15'd27349: duty=140; 15'd27350: duty=134; 15'd27351: duty=142;
15'd27352: duty=149; 15'd27353: duty=145; 15'd27354: duty=155; 15'd27355: duty=148; 15'd27356: duty=149; 15'd27357: duty=144; 15'd27358: duty=139; 15'd27359: duty=149;
15'd27360: duty=151; 15'd27361: duty=153; 15'd27362: duty=158; 15'd27363: duty=159; 15'd27364: duty=150; 15'd27365: duty=150; 15'd27366: duty=163; 15'd27367: duty=155;
15'd27368: duty=152; 15'd27369: duty=152; 15'd27370: duty=163; 15'd27371: duty=160; 15'd27372: duty=149; 15'd27373: duty=146; 15'd27374: duty=144; 15'd27375: duty=145;
15'd27376: duty=138; 15'd27377: duty=133; 15'd27378: duty=138; 15'd27379: duty=139; 15'd27380: duty=134; 15'd27381: duty=138; 15'd27382: duty=138; 15'd27383: duty=131;
15'd27384: duty=130; 15'd27385: duty=128; 15'd27386: duty=128; 15'd27387: duty=120; 15'd27388: duty=120; 15'd27389: duty=106; 15'd27390: duty=100; 15'd27391: duty=106;
15'd27392: duty=100; 15'd27393: duty=106; 15'd27394: duty=108; 15'd27395: duty=106; 15'd27396: duty=103; 15'd27397: duty=108; 15'd27398: duty=101; 15'd27399: duty=92;
15'd27400: duty=93; 15'd27401: duty=98; 15'd27402: duty=111; 15'd27403: duty=111; 15'd27404: duty=104; 15'd27405: duty=104; 15'd27406: duty=106; 15'd27407: duty=110;
15'd27408: duty=114; 15'd27409: duty=124; 15'd27410: duty=125; 15'd27411: duty=121; 15'd27412: duty=116; 15'd27413: duty=126; 15'd27414: duty=125; 15'd27415: duty=118;
15'd27416: duty=121; 15'd27417: duty=124; 15'd27418: duty=129; 15'd27419: duty=131; 15'd27420: duty=147; 15'd27421: duty=159; 15'd27422: duty=155; 15'd27423: duty=151;
15'd27424: duty=148; 15'd27425: duty=157; 15'd27426: duty=159; 15'd27427: duty=162; 15'd27428: duty=155; 15'd27429: duty=149; 15'd27430: duty=151; 15'd27431: duty=140;
15'd27432: duty=150; 15'd27433: duty=145; 15'd27434: duty=145; 15'd27435: duty=141; 15'd27436: duty=147; 15'd27437: duty=157; 15'd27438: duty=168; 15'd27439: duty=170;
15'd27440: duty=160; 15'd27441: duty=165; 15'd27442: duty=167; 15'd27443: duty=167; 15'd27444: duty=163; 15'd27445: duty=168; 15'd27446: duty=166; 15'd27447: duty=159;
15'd27448: duty=148; 15'd27449: duty=150; 15'd27450: duty=144; 15'd27451: duty=134; 15'd27452: duty=131; 15'd27453: duty=121; 15'd27454: duty=119; 15'd27455: duty=124;
15'd27456: duty=122; 15'd27457: duty=119; 15'd27458: duty=124; 15'd27459: duty=121; 15'd27460: duty=108; 15'd27461: duty=110; 15'd27462: duty=102; 15'd27463: duty=101;
15'd27464: duty=117; 15'd27465: duty=113; 15'd27466: duty=110; 15'd27467: duty=115; 15'd27468: duty=110; 15'd27469: duty=101; 15'd27470: duty=104; 15'd27471: duty=109;
15'd27472: duty=101; 15'd27473: duty=96; 15'd27474: duty=90; 15'd27475: duty=97; 15'd27476: duty=101; 15'd27477: duty=99; 15'd27478: duty=95; 15'd27479: duty=91;
15'd27480: duty=101; 15'd27481: duty=103; 15'd27482: duty=106; 15'd27483: duty=110; 15'd27484: duty=121; 15'd27485: duty=125; 15'd27486: duty=124; 15'd27487: duty=114;
15'd27488: duty=123; 15'd27489: duty=120; 15'd27490: duty=114; 15'd27491: duty=119; 15'd27492: duty=122; 15'd27493: duty=131; 15'd27494: duty=136; 15'd27495: duty=146;
15'd27496: duty=152; 15'd27497: duty=159; 15'd27498: duty=155; 15'd27499: duty=157; 15'd27500: duty=150; 15'd27501: duty=137; 15'd27502: duty=136; 15'd27503: duty=140;
15'd27504: duty=146; 15'd27505: duty=152; 15'd27506: duty=151; 15'd27507: duty=152; 15'd27508: duty=160; 15'd27509: duty=154; 15'd27510: duty=162; 15'd27511: duty=164;
15'd27512: duty=171; 15'd27513: duty=173; 15'd27514: duty=165; 15'd27515: duty=160; 15'd27516: duty=151; 15'd27517: duty=159; 15'd27518: duty=154; 15'd27519: duty=161;
15'd27520: duty=163; 15'd27521: duty=161; 15'd27522: duty=159; 15'd27523: duty=146; 15'd27524: duty=148; 15'd27525: duty=147; 15'd27526: duty=139; 15'd27527: duty=137;
15'd27528: duty=135; 15'd27529: duty=143; 15'd27530: duty=142; 15'd27531: duty=141; 15'd27532: duty=126; 15'd27533: duty=109; 15'd27534: duty=114; 15'd27535: duty=120;
15'd27536: duty=120; 15'd27537: duty=111; 15'd27538: duty=112; 15'd27539: duty=115; 15'd27540: duty=117; 15'd27541: duty=111; 15'd27542: duty=112; 15'd27543: duty=109;
15'd27544: duty=105; 15'd27545: duty=97; 15'd27546: duty=92; 15'd27547: duty=86; 15'd27548: duty=95; 15'd27549: duty=103; 15'd27550: duty=104; 15'd27551: duty=103;
15'd27552: duty=100; 15'd27553: duty=103; 15'd27554: duty=97; 15'd27555: duty=104; 15'd27556: duty=113; 15'd27557: duty=112; 15'd27558: duty=111; 15'd27559: duty=113;
15'd27560: duty=118; 15'd27561: duty=119; 15'd27562: duty=128; 15'd27563: duty=128; 15'd27564: duty=125; 15'd27565: duty=127; 15'd27566: duty=122; 15'd27567: duty=130;
15'd27568: duty=129; 15'd27569: duty=139; 15'd27570: duty=139; 15'd27571: duty=134; 15'd27572: duty=140; 15'd27573: duty=139; 15'd27574: duty=149; 15'd27575: duty=142;
15'd27576: duty=143; 15'd27577: duty=144; 15'd27578: duty=142; 15'd27579: duty=150; 15'd27580: duty=154; 15'd27581: duty=162; 15'd27582: duty=160; 15'd27583: duty=157;
15'd27584: duty=157; 15'd27585: duty=152; 15'd27586: duty=156; 15'd27587: duty=156; 15'd27588: duty=157; 15'd27589: duty=154; 15'd27590: duty=151; 15'd27591: duty=145;
15'd27592: duty=157; 15'd27593: duty=156; 15'd27594: duty=148; 15'd27595: duty=148; 15'd27596: duty=148; 15'd27597: duty=156; 15'd27598: duty=145; 15'd27599: duty=151;
15'd27600: duty=143; 15'd27601: duty=137; 15'd27602: duty=138; 15'd27603: duty=133; 15'd27604: duty=132; 15'd27605: duty=137; 15'd27606: duty=132; 15'd27607: duty=114;
15'd27608: duty=113; 15'd27609: duty=119; 15'd27610: duty=121; 15'd27611: duty=126; 15'd27612: duty=124; 15'd27613: duty=128; 15'd27614: duty=118; 15'd27615: duty=106;
15'd27616: duty=106; 15'd27617: duty=101; 15'd27618: duty=96; 15'd27619: duty=104; 15'd27620: duty=114; 15'd27621: duty=110; 15'd27622: duty=124; 15'd27623: duty=108;
15'd27624: duty=121; 15'd27625: duty=119; 15'd27626: duty=99; 15'd27627: duty=101; 15'd27628: duty=98; 15'd27629: duty=96; 15'd27630: duty=98; 15'd27631: duty=108;
15'd27632: duty=104; 15'd27633: duty=105; 15'd27634: duty=108; 15'd27635: duty=115; 15'd27636: duty=124; 15'd27637: duty=121; 15'd27638: duty=116; 15'd27639: duty=118;
15'd27640: duty=115; 15'd27641: duty=136; 15'd27642: duty=135; 15'd27643: duty=128; 15'd27644: duty=125; 15'd27645: duty=130; 15'd27646: duty=129; 15'd27647: duty=131;
15'd27648: duty=133; 15'd27649: duty=142; 15'd27650: duty=152; 15'd27651: duty=151; 15'd27652: duty=160; 15'd27653: duty=155; 15'd27654: duty=158; 15'd27655: duty=147;
15'd27656: duty=152; 15'd27657: duty=158; 15'd27658: duty=162; 15'd27659: duty=166; 15'd27660: duty=163; 15'd27661: duty=164; 15'd27662: duty=166; 15'd27663: duty=158;
15'd27664: duty=160; 15'd27665: duty=162; 15'd27666: duty=163; 15'd27667: duty=156; 15'd27668: duty=158; 15'd27669: duty=164; 15'd27670: duty=151; 15'd27671: duty=144;
15'd27672: duty=138; 15'd27673: duty=142; 15'd27674: duty=144; 15'd27675: duty=141; 15'd27676: duty=141; 15'd27677: duty=122; 15'd27678: duty=116; 15'd27679: duty=118;
15'd27680: duty=114; 15'd27681: duty=128; 15'd27682: duty=123; 15'd27683: duty=130; 15'd27684: duty=117; 15'd27685: duty=114; 15'd27686: duty=106; 15'd27687: duty=109;
15'd27688: duty=108; 15'd27689: duty=107; 15'd27690: duty=116; 15'd27691: duty=101; 15'd27692: duty=99; 15'd27693: duty=91; 15'd27694: duty=97; 15'd27695: duty=99;
15'd27696: duty=103; 15'd27697: duty=106; 15'd27698: duty=111; 15'd27699: duty=110; 15'd27700: duty=117; 15'd27701: duty=123; 15'd27702: duty=116; 15'd27703: duty=119;
15'd27704: duty=116; 15'd27705: duty=124; 15'd27706: duty=122; 15'd27707: duty=121; 15'd27708: duty=116; 15'd27709: duty=105; 15'd27710: duty=116; 15'd27711: duty=119;
15'd27712: duty=133; 15'd27713: duty=133; 15'd27714: duty=133; 15'd27715: duty=142; 15'd27716: duty=137; 15'd27717: duty=137; 15'd27718: duty=137; 15'd27719: duty=147;
15'd27720: duty=137; 15'd27721: duty=134; 15'd27722: duty=134; 15'd27723: duty=140; 15'd27724: duty=144; 15'd27725: duty=137; 15'd27726: duty=139; 15'd27727: duty=138;
15'd27728: duty=139; 15'd27729: duty=146; 15'd27730: duty=155; 15'd27731: duty=160; 15'd27732: duty=167; 15'd27733: duty=163; 15'd27734: duty=170; 15'd27735: duty=171;
15'd27736: duty=170; 15'd27737: duty=170; 15'd27738: duty=167; 15'd27739: duty=166; 15'd27740: duty=156; 15'd27741: duty=152; 15'd27742: duty=152; 15'd27743: duty=148;
15'd27744: duty=139; 15'd27745: duty=137; 15'd27746: duty=139; 15'd27747: duty=135; 15'd27748: duty=132; 15'd27749: duty=132; 15'd27750: duty=129; 15'd27751: duty=143;
15'd27752: duty=133; 15'd27753: duty=128; 15'd27754: duty=129; 15'd27755: duty=129; 15'd27756: duty=117; 15'd27757: duty=112; 15'd27758: duty=115; 15'd27759: duty=114;
15'd27760: duty=112; 15'd27761: duty=105; 15'd27762: duty=111; 15'd27763: duty=111; 15'd27764: duty=112; 15'd27765: duty=115; 15'd27766: duty=111; 15'd27767: duty=105;
15'd27768: duty=104; 15'd27769: duty=96; 15'd27770: duty=100; 15'd27771: duty=100; 15'd27772: duty=101; 15'd27773: duty=98; 15'd27774: duty=107; 15'd27775: duty=114;
15'd27776: duty=109; 15'd27777: duty=109; 15'd27778: duty=118; 15'd27779: duty=123; 15'd27780: duty=114; 15'd27781: duty=117; 15'd27782: duty=118; 15'd27783: duty=124;
15'd27784: duty=118; 15'd27785: duty=117; 15'd27786: duty=130; 15'd27787: duty=125; 15'd27788: duty=128; 15'd27789: duty=134; 15'd27790: duty=136; 15'd27791: duty=139;
15'd27792: duty=131; 15'd27793: duty=125; 15'd27794: duty=124; 15'd27795: duty=131; 15'd27796: duty=131; 15'd27797: duty=142; 15'd27798: duty=147; 15'd27799: duty=151;
15'd27800: duty=159; 15'd27801: duty=154; 15'd27802: duty=157; 15'd27803: duty=148; 15'd27804: duty=163; 15'd27805: duty=170; 15'd27806: duty=163; 15'd27807: duty=162;
15'd27808: duty=160; 15'd27809: duty=161; 15'd27810: duty=159; 15'd27811: duty=156; 15'd27812: duty=157; 15'd27813: duty=165; 15'd27814: duty=162; 15'd27815: duty=159;
15'd27816: duty=159; 15'd27817: duty=156; 15'd27818: duty=149; 15'd27819: duty=148; 15'd27820: duty=148; 15'd27821: duty=137; 15'd27822: duty=128; 15'd27823: duty=130;
15'd27824: duty=134; 15'd27825: duty=127; 15'd27826: duty=129; 15'd27827: duty=121; 15'd27828: duty=121; 15'd27829: duty=111; 15'd27830: duty=110; 15'd27831: duty=119;
15'd27832: duty=104; 15'd27833: duty=113; 15'd27834: duty=118; 15'd27835: duty=110; 15'd27836: duty=115; 15'd27837: duty=116; 15'd27838: duty=109; 15'd27839: duty=104;
15'd27840: duty=101; 15'd27841: duty=102; 15'd27842: duty=110; 15'd27843: duty=100; 15'd27844: duty=89; 15'd27845: duty=97; 15'd27846: duty=95; 15'd27847: duty=106;
15'd27848: duty=106; 15'd27849: duty=102; 15'd27850: duty=111; 15'd27851: duty=114; 15'd27852: duty=118; 15'd27853: duty=122; 15'd27854: duty=126; 15'd27855: duty=128;
15'd27856: duty=125; 15'd27857: duty=121; 15'd27858: duty=122; 15'd27859: duty=129; 15'd27860: duty=129; 15'd27861: duty=129; 15'd27862: duty=132; 15'd27863: duty=133;
15'd27864: duty=150; 15'd27865: duty=153; 15'd27866: duty=137; 15'd27867: duty=132; 15'd27868: duty=132; 15'd27869: duty=130; 15'd27870: duty=130; 15'd27871: duty=131;
15'd27872: duty=134; 15'd27873: duty=144; 15'd27874: duty=139; 15'd27875: duty=146; 15'd27876: duty=155; 15'd27877: duty=158; 15'd27878: duty=155; 15'd27879: duty=151;
15'd27880: duty=162; 15'd27881: duty=158; 15'd27882: duty=163; 15'd27883: duty=160; 15'd27884: duty=167; 15'd27885: duty=166; 15'd27886: duty=155; 15'd27887: duty=171;
15'd27888: duty=168; 15'd27889: duty=152; 15'd27890: duty=144; 15'd27891: duty=146; 15'd27892: duty=145; 15'd27893: duty=141; 15'd27894: duty=150; 15'd27895: duty=142;
15'd27896: duty=126; 15'd27897: duty=129; 15'd27898: duty=133; 15'd27899: duty=139; 15'd27900: duty=133; 15'd27901: duty=134; 15'd27902: duty=141; 15'd27903: duty=128;
15'd27904: duty=119; 15'd27905: duty=128; 15'd27906: duty=134; 15'd27907: duty=107; 15'd27908: duty=88; 15'd27909: duty=90; 15'd27910: duty=109; 15'd27911: duty=119;
15'd27912: duty=110; 15'd27913: duty=104; 15'd27914: duty=99; 15'd27915: duty=93; 15'd27916: duty=84; 15'd27917: duty=94; 15'd27918: duty=101; 15'd27919: duty=99;
15'd27920: duty=92; 15'd27921: duty=99; 15'd27922: duty=118; 15'd27923: duty=116; 15'd27924: duty=110; 15'd27925: duty=110; 15'd27926: duty=109; 15'd27927: duty=112;
15'd27928: duty=109; 15'd27929: duty=116; 15'd27930: duty=116; 15'd27931: duty=112; 15'd27932: duty=120; 15'd27933: duty=124; 15'd27934: duty=136; 15'd27935: duty=129;
15'd27936: duty=128; 15'd27937: duty=131; 15'd27938: duty=142; 15'd27939: duty=159; 15'd27940: duty=153; 15'd27941: duty=152; 15'd27942: duty=148; 15'd27943: duty=140;
15'd27944: duty=142; 15'd27945: duty=137; 15'd27946: duty=140; 15'd27947: duty=157; 15'd27948: duty=154; 15'd27949: duty=156; 15'd27950: duty=162; 15'd27951: duty=153;
15'd27952: duty=161; 15'd27953: duty=160; 15'd27954: duty=149; 15'd27955: duty=157; 15'd27956: duty=159; 15'd27957: duty=159; 15'd27958: duty=165; 15'd27959: duty=154;
15'd27960: duty=156; 15'd27961: duty=160; 15'd27962: duty=160; 15'd27963: duty=157; 15'd27964: duty=159; 15'd27965: duty=159; 15'd27966: duty=156; 15'd27967: duty=151;
15'd27968: duty=145; 15'd27969: duty=147; 15'd27970: duty=124; 15'd27971: duty=119; 15'd27972: duty=110; 15'd27973: duty=118; 15'd27974: duty=118; 15'd27975: duty=121;
15'd27976: duty=125; 15'd27977: duty=112; 15'd27978: duty=119; 15'd27979: duty=113; 15'd27980: duty=125; 15'd27981: duty=127; 15'd27982: duty=115; 15'd27983: duty=105;
15'd27984: duty=110; 15'd27985: duty=107; 15'd27986: duty=85; 15'd27987: duty=85; 15'd27988: duty=91; 15'd27989: duty=99; 15'd27990: duty=98; 15'd27991: duty=98;
15'd27992: duty=107; 15'd27993: duty=108; 15'd27994: duty=114; 15'd27995: duty=109; 15'd27996: duty=112; 15'd27997: duty=113; 15'd27998: duty=110; 15'd27999: duty=110;
15'd28000: duty=113; 15'd28001: duty=112; 15'd28002: duty=108; 15'd28003: duty=104; 15'd28004: duty=105; 15'd28005: duty=118; 15'd28006: duty=111; 15'd28007: duty=125;
15'd28008: duty=128; 15'd28009: duty=128; 15'd28010: duty=145; 15'd28011: duty=140; 15'd28012: duty=140; 15'd28013: duty=134; 15'd28014: duty=124; 15'd28015: duty=137;
15'd28016: duty=140; 15'd28017: duty=134; 15'd28018: duty=146; 15'd28019: duty=148; 15'd28020: duty=143; 15'd28021: duty=139; 15'd28022: duty=142; 15'd28023: duty=154;
15'd28024: duty=163; 15'd28025: duty=168; 15'd28026: duty=172; 15'd28027: duty=176; 15'd28028: duty=171; 15'd28029: duty=169; 15'd28030: duty=168; 15'd28031: duty=164;
15'd28032: duty=157; 15'd28033: duty=159; 15'd28034: duty=160; 15'd28035: duty=152; 15'd28036: duty=152; 15'd28037: duty=141; 15'd28038: duty=154; 15'd28039: duty=149;
15'd28040: duty=154; 15'd28041: duty=161; 15'd28042: duty=150; 15'd28043: duty=150; 15'd28044: duty=137; 15'd28045: duty=136; 15'd28046: duty=122; 15'd28047: duty=121;
15'd28048: duty=113; 15'd28049: duty=125; 15'd28050: duty=134; 15'd28051: duty=123; 15'd28052: duty=126; 15'd28053: duty=118; 15'd28054: duty=120; 15'd28055: duty=130;
15'd28056: duty=120; 15'd28057: duty=117; 15'd28058: duty=123; 15'd28059: duty=107; 15'd28060: duty=111; 15'd28061: duty=112; 15'd28062: duty=99; 15'd28063: duty=97;
15'd28064: duty=97; 15'd28065: duty=98; 15'd28066: duty=101; 15'd28067: duty=101; 15'd28068: duty=94; 15'd28069: duty=101; 15'd28070: duty=99; 15'd28071: duty=93;
15'd28072: duty=105; 15'd28073: duty=103; 15'd28074: duty=107; 15'd28075: duty=124; 15'd28076: duty=108; 15'd28077: duty=99; 15'd28078: duty=110; 15'd28079: duty=106;
15'd28080: duty=110; 15'd28081: duty=118; 15'd28082: duty=121; 15'd28083: duty=126; 15'd28084: duty=131; 15'd28085: duty=127; 15'd28086: duty=128; 15'd28087: duty=132;
15'd28088: duty=132; 15'd28089: duty=147; 15'd28090: duty=151; 15'd28091: duty=150; 15'd28092: duty=152; 15'd28093: duty=145; 15'd28094: duty=148; 15'd28095: duty=158;
15'd28096: duty=162; 15'd28097: duty=162; 15'd28098: duty=169; 15'd28099: duty=166; 15'd28100: duty=165; 15'd28101: duty=164; 15'd28102: duty=155; 15'd28103: duty=168;
15'd28104: duty=166; 15'd28105: duty=164; 15'd28106: duty=169; 15'd28107: duty=164; 15'd28108: duty=158; 15'd28109: duty=152; 15'd28110: duty=141; 15'd28111: duty=155;
15'd28112: duty=155; 15'd28113: duty=143; 15'd28114: duty=137; 15'd28115: duty=129; 15'd28116: duty=135; 15'd28117: duty=130; 15'd28118: duty=115; 15'd28119: duty=118;
15'd28120: duty=123; 15'd28121: duty=116; 15'd28122: duty=117; 15'd28123: duty=123; 15'd28124: duty=119; 15'd28125: duty=123; 15'd28126: duty=126; 15'd28127: duty=122;
15'd28128: duty=123; 15'd28129: duty=117; 15'd28130: duty=118; 15'd28131: duty=104; 15'd28132: duty=96; 15'd28133: duty=87; 15'd28134: duty=103; 15'd28135: duty=112;
15'd28136: duty=94; 15'd28137: duty=101; 15'd28138: duty=111; 15'd28139: duty=114; 15'd28140: duty=111; 15'd28141: duty=107; 15'd28142: duty=110; 15'd28143: duty=121;
15'd28144: duty=126; 15'd28145: duty=128; 15'd28146: duty=120; 15'd28147: duty=110; 15'd28148: duty=111; 15'd28149: duty=107; 15'd28150: duty=117; 15'd28151: duty=136;
15'd28152: duty=129; 15'd28153: duty=133; 15'd28154: duty=136; 15'd28155: duty=135; 15'd28156: duty=139; 15'd28157: duty=136; 15'd28158: duty=142; 15'd28159: duty=155;
15'd28160: duty=155; 15'd28161: duty=142; 15'd28162: duty=145; 15'd28163: duty=135; 15'd28164: duty=129; 15'd28165: duty=130; 15'd28166: duty=130; 15'd28167: duty=142;
15'd28168: duty=143; 15'd28169: duty=142; 15'd28170: duty=147; 15'd28171: duty=154; 15'd28172: duty=153; 15'd28173: duty=164; 15'd28174: duty=157; 15'd28175: duty=154;
15'd28176: duty=154; 15'd28177: duty=157; 15'd28178: duty=148; 15'd28179: duty=155; 15'd28180: duty=153; 15'd28181: duty=142; 15'd28182: duty=145; 15'd28183: duty=131;
15'd28184: duty=128; 15'd28185: duty=140; 15'd28186: duty=141; 15'd28187: duty=128; 15'd28188: duty=144; 15'd28189: duty=124; 15'd28190: duty=126; 15'd28191: duty=127;
15'd28192: duty=134; 15'd28193: duty=139; 15'd28194: duty=138; 15'd28195: duty=135; 15'd28196: duty=126; 15'd28197: duty=131; 15'd28198: duty=131; 15'd28199: duty=134;
15'd28200: duty=126; 15'd28201: duty=131; 15'd28202: duty=127; 15'd28203: duty=118; 15'd28204: duty=105; 15'd28205: duty=119; 15'd28206: duty=113; 15'd28207: duty=102;
15'd28208: duty=102; 15'd28209: duty=102; 15'd28210: duty=115; 15'd28211: duty=102; 15'd28212: duty=106; 15'd28213: duty=110; 15'd28214: duty=110; 15'd28215: duty=122;
15'd28216: duty=123; 15'd28217: duty=111; 15'd28218: duty=110; 15'd28219: duty=113; 15'd28220: duty=116; 15'd28221: duty=124; 15'd28222: duty=122; 15'd28223: duty=122;
15'd28224: duty=116; 15'd28225: duty=124; 15'd28226: duty=118; 15'd28227: duty=125; 15'd28228: duty=134; 15'd28229: duty=129; 15'd28230: duty=134; 15'd28231: duty=122;
15'd28232: duty=124; 15'd28233: duty=120; 15'd28234: duty=121; 15'd28235: duty=137; 15'd28236: duty=133; 15'd28237: duty=131; 15'd28238: duty=145; 15'd28239: duty=148;
15'd28240: duty=150; 15'd28241: duty=154; 15'd28242: duty=156; 15'd28243: duty=151; 15'd28244: duty=152; 15'd28245: duty=156; 15'd28246: duty=159; 15'd28247: duty=159;
15'd28248: duty=150; 15'd28249: duty=154; 15'd28250: duty=154; 15'd28251: duty=149; 15'd28252: duty=154; 15'd28253: duty=149; 15'd28254: duty=145; 15'd28255: duty=147;
15'd28256: duty=139; 15'd28257: duty=145; 15'd28258: duty=147; 15'd28259: duty=142; 15'd28260: duty=147; 15'd28261: duty=143; 15'd28262: duty=138; 15'd28263: duty=129;
15'd28264: duty=134; 15'd28265: duty=137; 15'd28266: duty=124; 15'd28267: duty=124; 15'd28268: duty=124; 15'd28269: duty=125; 15'd28270: duty=126; 15'd28271: duty=112;
15'd28272: duty=118; 15'd28273: duty=124; 15'd28274: duty=119; 15'd28275: duty=128; 15'd28276: duty=131; 15'd28277: duty=131; 15'd28278: duty=131; 15'd28279: duty=120;
15'd28280: duty=102; 15'd28281: duty=105; 15'd28282: duty=99; 15'd28283: duty=113; 15'd28284: duty=118; 15'd28285: duty=109; 15'd28286: duty=115; 15'd28287: duty=110;
15'd28288: duty=116; 15'd28289: duty=113; 15'd28290: duty=115; 15'd28291: duty=118; 15'd28292: duty=113; 15'd28293: duty=112; 15'd28294: duty=119; 15'd28295: duty=116;
15'd28296: duty=119; 15'd28297: duty=120; 15'd28298: duty=118; 15'd28299: duty=124; 15'd28300: duty=127; 15'd28301: duty=128; 15'd28302: duty=134; 15'd28303: duty=139;
15'd28304: duty=136; 15'd28305: duty=145; 15'd28306: duty=134; 15'd28307: duty=134; 15'd28308: duty=128; 15'd28309: duty=128; 15'd28310: duty=134; 15'd28311: duty=128;
15'd28312: duty=129; 15'd28313: duty=134; 15'd28314: duty=139; 15'd28315: duty=145; 15'd28316: duty=142; 15'd28317: duty=149; 15'd28318: duty=157; 15'd28319: duty=156;
15'd28320: duty=160; 15'd28321: duty=153; 15'd28322: duty=149; 15'd28323: duty=153; 15'd28324: duty=160; 15'd28325: duty=148; 15'd28326: duty=151; 15'd28327: duty=153;
15'd28328: duty=151; 15'd28329: duty=151; 15'd28330: duty=142; 15'd28331: duty=138; 15'd28332: duty=139; 15'd28333: duty=137; 15'd28334: duty=136; 15'd28335: duty=137;
15'd28336: duty=131; 15'd28337: duty=127; 15'd28338: duty=128; 15'd28339: duty=114; 15'd28340: duty=120; 15'd28341: duty=110; 15'd28342: duty=114; 15'd28343: duty=118;
15'd28344: duty=111; 15'd28345: duty=127; 15'd28346: duty=137; 15'd28347: duty=142; 15'd28348: duty=122; 15'd28349: duty=124; 15'd28350: duty=122; 15'd28351: duty=118;
15'd28352: duty=113; 15'd28353: duty=106; 15'd28354: duty=102; 15'd28355: duty=108; 15'd28356: duty=115; 15'd28357: duty=115; 15'd28358: duty=115; 15'd28359: duty=115;
15'd28360: duty=106; 15'd28361: duty=112; 15'd28362: duty=104; 15'd28363: duty=110; 15'd28364: duty=127; 15'd28365: duty=119; 15'd28366: duty=119; 15'd28367: duty=115;
15'd28368: duty=116; 15'd28369: duty=113; 15'd28370: duty=118; 15'd28371: duty=125; 15'd28372: duty=126; 15'd28373: duty=134; 15'd28374: duty=136; 15'd28375: duty=134;
15'd28376: duty=131; 15'd28377: duty=131; 15'd28378: duty=131; 15'd28379: duty=130; 15'd28380: duty=139; 15'd28381: duty=148; 15'd28382: duty=155; 15'd28383: duty=148;
15'd28384: duty=151; 15'd28385: duty=153; 15'd28386: duty=149; 15'd28387: duty=157; 15'd28388: duty=165; 15'd28389: duty=168; 15'd28390: duty=163; 15'd28391: duty=162;
15'd28392: duty=165; 15'd28393: duty=171; 15'd28394: duty=167; 15'd28395: duty=165; 15'd28396: duty=162; 15'd28397: duty=161; 15'd28398: duty=163; 15'd28399: duty=153;
15'd28400: duty=160; 15'd28401: duty=161; 15'd28402: duty=149; 15'd28403: duty=135; 15'd28404: duty=125; 15'd28405: duty=126; 15'd28406: duty=130; 15'd28407: duty=124;
15'd28408: duty=117; 15'd28409: duty=115; 15'd28410: duty=117; 15'd28411: duty=110; 15'd28412: duty=106; 15'd28413: duty=104; 15'd28414: duty=108; 15'd28415: duty=112;
15'd28416: duty=104; 15'd28417: duty=120; 15'd28418: duty=102; 15'd28419: duty=106; 15'd28420: duty=97; 15'd28421: duty=90; 15'd28422: duty=100; 15'd28423: duty=95;
15'd28424: duty=96; 15'd28425: duty=89; 15'd28426: duty=90; 15'd28427: duty=90; 15'd28428: duty=93; 15'd28429: duty=97; 15'd28430: duty=110; 15'd28431: duty=102;
15'd28432: duty=104; 15'd28433: duty=121; 15'd28434: duty=107; 15'd28435: duty=113; 15'd28436: duty=116; 15'd28437: duty=104; 15'd28438: duty=118; 15'd28439: duty=122;
15'd28440: duty=119; 15'd28441: duty=121; 15'd28442: duty=121; 15'd28443: duty=142; 15'd28444: duty=147; 15'd28445: duty=148; 15'd28446: duty=153; 15'd28447: duty=149;
15'd28448: duty=147; 15'd28449: duty=146; 15'd28450: duty=148; 15'd28451: duty=149; 15'd28452: duty=148; 15'd28453: duty=135; 15'd28454: duty=139; 15'd28455: duty=143;
15'd28456: duty=151; 15'd28457: duty=151; 15'd28458: duty=161; 15'd28459: duty=157; 15'd28460: duty=167; 15'd28461: duty=171; 15'd28462: duty=176; 15'd28463: duty=185;
15'd28464: duty=179; 15'd28465: duty=162; 15'd28466: duty=162; 15'd28467: duty=165; 15'd28468: duty=163; 15'd28469: duty=172; 15'd28470: duty=159; 15'd28471: duty=157;
15'd28472: duty=154; 15'd28473: duty=151; 15'd28474: duty=153; 15'd28475: duty=165; 15'd28476: duty=153; 15'd28477: duty=156; 15'd28478: duty=139; 15'd28479: duty=141;
15'd28480: duty=148; 15'd28481: duty=140; 15'd28482: duty=128; 15'd28483: duty=114; 15'd28484: duty=116; 15'd28485: duty=116; 15'd28486: duty=113; 15'd28487: duty=96;
15'd28488: duty=111; 15'd28489: duty=118; 15'd28490: duty=111; 15'd28491: duty=114; 15'd28492: duty=105; 15'd28493: duty=99; 15'd28494: duty=109; 15'd28495: duty=92;
15'd28496: duty=91; 15'd28497: duty=92; 15'd28498: duty=89; 15'd28499: duty=104; 15'd28500: duty=94; 15'd28501: duty=101; 15'd28502: duty=99; 15'd28503: duty=93;
15'd28504: duty=90; 15'd28505: duty=102; 15'd28506: duty=105; 15'd28507: duty=99; 15'd28508: duty=104; 15'd28509: duty=109; 15'd28510: duty=115; 15'd28511: duty=112;
15'd28512: duty=113; 15'd28513: duty=115; 15'd28514: duty=126; 15'd28515: duty=133; 15'd28516: duty=136; 15'd28517: duty=145; 15'd28518: duty=149; 15'd28519: duty=133;
15'd28520: duty=143; 15'd28521: duty=137; 15'd28522: duty=134; 15'd28523: duty=129; 15'd28524: duty=127; 15'd28525: duty=137; 15'd28526: duty=136; 15'd28527: duty=136;
15'd28528: duty=148; 15'd28529: duty=149; 15'd28530: duty=159; 15'd28531: duty=163; 15'd28532: duty=159; 15'd28533: duty=174; 15'd28534: duty=173; 15'd28535: duty=173;
15'd28536: duty=160; 15'd28537: duty=162; 15'd28538: duty=151; 15'd28539: duty=155; 15'd28540: duty=157; 15'd28541: duty=159; 15'd28542: duty=156; 15'd28543: duty=145;
15'd28544: duty=148; 15'd28545: duty=156; 15'd28546: duty=151; 15'd28547: duty=151; 15'd28548: duty=149; 15'd28549: duty=142; 15'd28550: duty=140; 15'd28551: duty=137;
15'd28552: duty=145; 15'd28553: duty=144; 15'd28554: duty=121; 15'd28555: duty=104; 15'd28556: duty=105; 15'd28557: duty=113; 15'd28558: duty=122; 15'd28559: duty=110;
15'd28560: duty=107; 15'd28561: duty=107; 15'd28562: duty=115; 15'd28563: duty=115; 15'd28564: duty=111; 15'd28565: duty=118; 15'd28566: duty=115; 15'd28567: duty=92;
15'd28568: duty=96; 15'd28569: duty=104; 15'd28570: duty=92; 15'd28571: duty=96; 15'd28572: duty=100; 15'd28573: duty=105; 15'd28574: duty=110; 15'd28575: duty=113;
15'd28576: duty=106; 15'd28577: duty=111; 15'd28578: duty=115; 15'd28579: duty=116; 15'd28580: duty=124; 15'd28581: duty=125; 15'd28582: duty=131; 15'd28583: duty=134;
15'd28584: duty=128; 15'd28585: duty=124; 15'd28586: duty=120; 15'd28587: duty=120; 15'd28588: duty=124; 15'd28589: duty=128; 15'd28590: duty=147; 15'd28591: duty=147;
15'd28592: duty=149; 15'd28593: duty=154; 15'd28594: duty=156; 15'd28595: duty=157; 15'd28596: duty=147; 15'd28597: duty=149; 15'd28598: duty=150; 15'd28599: duty=137;
15'd28600: duty=141; 15'd28601: duty=140; 15'd28602: duty=141; 15'd28603: duty=146; 15'd28604: duty=145; 15'd28605: duty=154; 15'd28606: duty=155; 15'd28607: duty=161;
15'd28608: duty=158; 15'd28609: duty=167; 15'd28610: duty=171; 15'd28611: duty=166; 15'd28612: duty=155; 15'd28613: duty=151; 15'd28614: duty=147; 15'd28615: duty=141;
15'd28616: duty=147; 15'd28617: duty=149; 15'd28618: duty=142; 15'd28619: duty=152; 15'd28620: duty=145; 15'd28621: duty=137; 15'd28622: duty=140; 15'd28623: duty=130;
15'd28624: duty=135; 15'd28625: duty=122; 15'd28626: duty=137; 15'd28627: duty=129; 15'd28628: duty=117; 15'd28629: duty=102; 15'd28630: duty=99; 15'd28631: duty=108;
15'd28632: duty=107; 15'd28633: duty=124; 15'd28634: duty=120; 15'd28635: duty=119; 15'd28636: duty=114; 15'd28637: duty=112; 15'd28638: duty=113; 15'd28639: duty=110;
15'd28640: duty=111; 15'd28641: duty=121; 15'd28642: duty=110; 15'd28643: duty=101; 15'd28644: duty=105; 15'd28645: duty=96; 15'd28646: duty=96; 15'd28647: duty=96;
15'd28648: duty=99; 15'd28649: duty=101; 15'd28650: duty=99; 15'd28651: duty=110; 15'd28652: duty=116; 15'd28653: duty=121; 15'd28654: duty=121; 15'd28655: duty=117;
15'd28656: duty=117; 15'd28657: duty=127; 15'd28658: duty=126; 15'd28659: duty=114; 15'd28660: duty=124; 15'd28661: duty=121; 15'd28662: duty=128; 15'd28663: duty=130;
15'd28664: duty=136; 15'd28665: duty=149; 15'd28666: duty=145; 15'd28667: duty=138; 15'd28668: duty=135; 15'd28669: duty=133; 15'd28670: duty=131; 15'd28671: duty=133;
15'd28672: duty=131; 15'd28673: duty=132; 15'd28674: duty=136; 15'd28675: duty=148; 15'd28676: duty=164; 15'd28677: duty=162; 15'd28678: duty=169; 15'd28679: duty=179;
15'd28680: duty=177; 15'd28681: duty=159; 15'd28682: duty=156; 15'd28683: duty=152; 15'd28684: duty=151; 15'd28685: duty=160; 15'd28686: duty=157; 15'd28687: duty=168;
15'd28688: duty=157; 15'd28689: duty=154; 15'd28690: duty=154; 15'd28691: duty=162; 15'd28692: duty=162; 15'd28693: duty=151; 15'd28694: duty=142; 15'd28695: duty=145;
15'd28696: duty=145; 15'd28697: duty=142; 15'd28698: duty=147; 15'd28699: duty=132; 15'd28700: duty=124; 15'd28701: duty=114; 15'd28702: duty=119; 15'd28703: duty=126;
15'd28704: duty=118; 15'd28705: duty=114; 15'd28706: duty=127; 15'd28707: duty=125; 15'd28708: duty=116; 15'd28709: duty=113; 15'd28710: duty=115; 15'd28711: duty=123;
15'd28712: duty=115; 15'd28713: duty=105; 15'd28714: duty=107; 15'd28715: duty=99; 15'd28716: duty=79; 15'd28717: duty=93; 15'd28718: duty=82; 15'd28719: duty=91;
15'd28720: duty=102; 15'd28721: duty=96; 15'd28722: duty=104; 15'd28723: duty=113; 15'd28724: duty=110; 15'd28725: duty=113; 15'd28726: duty=116; 15'd28727: duty=111;
15'd28728: duty=120; 15'd28729: duty=120; 15'd28730: duty=121; 15'd28731: duty=118; 15'd28732: duty=123; 15'd28733: duty=129; 15'd28734: duty=126; 15'd28735: duty=137;
15'd28736: duty=148; 15'd28737: duty=148; 15'd28738: duty=142; 15'd28739: duty=143; 15'd28740: duty=145; 15'd28741: duty=134; 15'd28742: duty=132; 15'd28743: duty=135;
15'd28744: duty=134; 15'd28745: duty=132; 15'd28746: duty=136; 15'd28747: duty=143; 15'd28748: duty=145; 15'd28749: duty=148; 15'd28750: duty=159; 15'd28751: duty=160;
15'd28752: duty=170; 15'd28753: duty=168; 15'd28754: duty=155; 15'd28755: duty=159; 15'd28756: duty=148; 15'd28757: duty=144; 15'd28758: duty=160; 15'd28759: duty=150;
15'd28760: duty=151; 15'd28761: duty=154; 15'd28762: duty=148; 15'd28763: duty=148; 15'd28764: duty=140; 15'd28765: duty=144; 15'd28766: duty=145; 15'd28767: duty=142;
15'd28768: duty=131; 15'd28769: duty=131; 15'd28770: duty=122; 15'd28771: duty=124; 15'd28772: duty=116; 15'd28773: duty=123; 15'd28774: duty=128; 15'd28775: duty=130;
15'd28776: duty=125; 15'd28777: duty=118; 15'd28778: duty=131; 15'd28779: duty=125; 15'd28780: duty=141; 15'd28781: duty=124; 15'd28782: duty=109; 15'd28783: duty=113;
15'd28784: duty=114; 15'd28785: duty=109; 15'd28786: duty=109; 15'd28787: duty=101; 15'd28788: duty=91; 15'd28789: duty=95; 15'd28790: duty=90; 15'd28791: duty=105;
15'd28792: duty=106; 15'd28793: duty=108; 15'd28794: duty=114; 15'd28795: duty=114; 15'd28796: duty=112; 15'd28797: duty=109; 15'd28798: duty=116; 15'd28799: duty=117;
15'd28800: duty=125; 15'd28801: duty=126; 15'd28802: duty=129; 15'd28803: duty=115; 15'd28804: duty=123; 15'd28805: duty=133; 15'd28806: duty=138; 15'd28807: duty=142;
15'd28808: duty=132; 15'd28809: duty=147; 15'd28810: duty=139; 15'd28811: duty=144; 15'd28812: duty=151; 15'd28813: duty=148; 15'd28814: duty=134; 15'd28815: duty=134;
15'd28816: duty=134; 15'd28817: duty=136; 15'd28818: duty=146; 15'd28819: duty=142; 15'd28820: duty=153; 15'd28821: duty=153; 15'd28822: duty=159; 15'd28823: duty=160;
15'd28824: duty=169; 15'd28825: duty=167; 15'd28826: duty=153; 15'd28827: duty=162; 15'd28828: duty=165; 15'd28829: duty=160; 15'd28830: duty=148; 15'd28831: duty=147;
15'd28832: duty=142; 15'd28833: duty=140; 15'd28834: duty=141; 15'd28835: duty=140; 15'd28836: duty=140; 15'd28837: duty=145; 15'd28838: duty=153; 15'd28839: duty=147;
15'd28840: duty=133; 15'd28841: duty=125; 15'd28842: duty=122; 15'd28843: duty=119; 15'd28844: duty=119; 15'd28845: duty=109; 15'd28846: duty=117; 15'd28847: duty=116;
15'd28848: duty=113; 15'd28849: duty=112; 15'd28850: duty=113; 15'd28851: duty=116; 15'd28852: duty=114; 15'd28853: duty=106; 15'd28854: duty=105; 15'd28855: duty=116;
15'd28856: duty=109; 15'd28857: duty=107; 15'd28858: duty=99; 15'd28859: duty=103; 15'd28860: duty=104; 15'd28861: duty=106; 15'd28862: duty=106; 15'd28863: duty=96;
15'd28864: duty=108; 15'd28865: duty=101; 15'd28866: duty=105; 15'd28867: duty=108; 15'd28868: duty=108; 15'd28869: duty=118; 15'd28870: duty=112; 15'd28871: duty=122;
15'd28872: duty=133; 15'd28873: duty=133; 15'd28874: duty=117; 15'd28875: duty=103; 15'd28876: duty=110; 15'd28877: duty=122; 15'd28878: duty=132; 15'd28879: duty=141;
15'd28880: duty=144; 15'd28881: duty=146; 15'd28882: duty=147; 15'd28883: duty=142; 15'd28884: duty=138; 15'd28885: duty=151; 15'd28886: duty=141; 15'd28887: duty=131;
15'd28888: duty=137; 15'd28889: duty=133; 15'd28890: duty=145; 15'd28891: duty=142; 15'd28892: duty=140; 15'd28893: duty=157; 15'd28894: duty=162; 15'd28895: duty=156;
15'd28896: duty=162; 15'd28897: duty=165; 15'd28898: duty=163; 15'd28899: duty=166; 15'd28900: duty=167; 15'd28901: duty=154; 15'd28902: duty=150; 15'd28903: duty=146;
15'd28904: duty=152; 15'd28905: duty=152; 15'd28906: duty=156; 15'd28907: duty=151; 15'd28908: duty=150; 15'd28909: duty=158; 15'd28910: duty=153; 15'd28911: duty=151;
15'd28912: duty=130; 15'd28913: duty=140; 15'd28914: duty=135; 15'd28915: duty=127; 15'd28916: duty=132; 15'd28917: duty=128; 15'd28918: duty=124; 15'd28919: duty=116;
15'd28920: duty=100; 15'd28921: duty=107; 15'd28922: duty=126; 15'd28923: duty=114; 15'd28924: duty=125; 15'd28925: duty=134; 15'd28926: duty=121; 15'd28927: duty=134;
15'd28928: duty=128; 15'd28929: duty=121; 15'd28930: duty=128; 15'd28931: duty=121; 15'd28932: duty=119; 15'd28933: duty=114; 15'd28934: duty=100; 15'd28935: duty=98;
15'd28936: duty=105; 15'd28937: duty=113; 15'd28938: duty=115; 15'd28939: duty=104; 15'd28940: duty=107; 15'd28941: duty=109; 15'd28942: duty=105; 15'd28943: duty=102;
15'd28944: duty=102; 15'd28945: duty=108; 15'd28946: duty=115; 15'd28947: duty=118; 15'd28948: duty=113; 15'd28949: duty=116; 15'd28950: duty=124; 15'd28951: duty=124;
15'd28952: duty=121; 15'd28953: duty=123; 15'd28954: duty=132; 15'd28955: duty=133; 15'd28956: duty=129; 15'd28957: duty=118; 15'd28958: duty=124; 15'd28959: duty=127;
15'd28960: duty=122; 15'd28961: duty=124; 15'd28962: duty=128; 15'd28963: duty=128; 15'd28964: duty=138; 15'd28965: duty=148; 15'd28966: duty=144; 15'd28967: duty=153;
15'd28968: duty=159; 15'd28969: duty=164; 15'd28970: duty=164; 15'd28971: duty=166; 15'd28972: duty=160; 15'd28973: duty=162; 15'd28974: duty=162; 15'd28975: duty=161;
15'd28976: duty=159; 15'd28977: duty=163; 15'd28978: duty=158; 15'd28979: duty=143; 15'd28980: duty=136; 15'd28981: duty=154; 15'd28982: duty=165; 15'd28983: duty=153;
15'd28984: duty=148; 15'd28985: duty=136; 15'd28986: duty=135; 15'd28987: duty=133; 15'd28988: duty=136; 15'd28989: duty=133; 15'd28990: duty=125; 15'd28991: duty=117;
15'd28992: duty=113; 15'd28993: duty=124; 15'd28994: duty=127; 15'd28995: duty=122; 15'd28996: duty=118; 15'd28997: duty=106; 15'd28998: duty=112; 15'd28999: duty=118;
15'd29000: duty=131; 15'd29001: duty=127; 15'd29002: duty=108; 15'd29003: duty=104; 15'd29004: duty=102; 15'd29005: duty=118; 15'd29006: duty=107; 15'd29007: duty=97;
15'd29008: duty=110; 15'd29009: duty=116; 15'd29010: duty=124; 15'd29011: duty=121; 15'd29012: duty=122; 15'd29013: duty=113; 15'd29014: duty=116; 15'd29015: duty=110;
15'd29016: duty=104; 15'd29017: duty=115; 15'd29018: duty=113; 15'd29019: duty=127; 15'd29020: duty=122; 15'd29021: duty=124; 15'd29022: duty=119; 15'd29023: duty=124;
15'd29024: duty=134; 15'd29025: duty=142; 15'd29026: duty=143; 15'd29027: duty=137; 15'd29028: duty=155; 15'd29029: duty=140; 15'd29030: duty=134; 15'd29031: duty=127;
15'd29032: duty=113; 15'd29033: duty=127; 15'd29034: duty=127; 15'd29035: duty=133; 15'd29036: duty=139; 15'd29037: duty=134; 15'd29038: duty=138; 15'd29039: duty=140;
15'd29040: duty=146; 15'd29041: duty=152; 15'd29042: duty=165; 15'd29043: duty=164; 15'd29044: duty=166; 15'd29045: duty=156; 15'd29046: duty=142; 15'd29047: duty=151;
15'd29048: duty=150; 15'd29049: duty=153; 15'd29050: duty=156; 15'd29051: duty=152; 15'd29052: duty=147; 15'd29053: duty=148; 15'd29054: duty=151; 15'd29055: duty=151;
15'd29056: duty=151; 15'd29057: duty=148; 15'd29058: duty=147; 15'd29059: duty=145; 15'd29060: duty=136; 15'd29061: duty=129; 15'd29062: duty=119; 15'd29063: duty=127;
15'd29064: duty=133; 15'd29065: duty=124; 15'd29066: duty=126; 15'd29067: duty=137; 15'd29068: duty=131; 15'd29069: duty=129; 15'd29070: duty=130; 15'd29071: duty=121;
15'd29072: duty=123; 15'd29073: duty=113; 15'd29074: duty=99; 15'd29075: duty=102; 15'd29076: duty=103; 15'd29077: duty=94; 15'd29078: duty=95; 15'd29079: duty=81;
15'd29080: duty=98; 15'd29081: duty=101; 15'd29082: duty=98; 15'd29083: duty=112; 15'd29084: duty=104; 15'd29085: duty=104; 15'd29086: duty=107; 15'd29087: duty=108;
15'd29088: duty=110; 15'd29089: duty=115; 15'd29090: duty=107; 15'd29091: duty=115; 15'd29092: duty=111; 15'd29093: duty=114; 15'd29094: duty=121; 15'd29095: duty=124;
15'd29096: duty=121; 15'd29097: duty=114; 15'd29098: duty=116; 15'd29099: duty=133; 15'd29100: duty=137; 15'd29101: duty=123; 15'd29102: duty=131; 15'd29103: duty=127;
15'd29104: duty=131; 15'd29105: duty=135; 15'd29106: duty=132; 15'd29107: duty=155; 15'd29108: duty=151; 15'd29109: duty=155; 15'd29110: duty=160; 15'd29111: duty=148;
15'd29112: duty=156; 15'd29113: duty=161; 15'd29114: duty=165; 15'd29115: duty=164; 15'd29116: duty=164; 15'd29117: duty=173; 15'd29118: duty=184; 15'd29119: duty=170;
15'd29120: duty=171; 15'd29121: duty=154; 15'd29122: duty=154; 15'd29123: duty=170; 15'd29124: duty=171; 15'd29125: duty=163; 15'd29126: duty=153; 15'd29127: duty=151;
15'd29128: duty=150; 15'd29129: duty=151; 15'd29130: duty=130; 15'd29131: duty=126; 15'd29132: duty=128; 15'd29133: duty=135; 15'd29134: duty=142; 15'd29135: duty=132;
15'd29136: duty=113; 15'd29137: duty=117; 15'd29138: duty=129; 15'd29139: duty=127; 15'd29140: duty=122; 15'd29141: duty=122; 15'd29142: duty=110; 15'd29143: duty=108;
15'd29144: duty=114; 15'd29145: duty=119; 15'd29146: duty=130; 15'd29147: duty=114; 15'd29148: duty=100; 15'd29149: duty=106; 15'd29150: duty=104; 15'd29151: duty=96;
15'd29152: duty=88; 15'd29153: duty=90; 15'd29154: duty=93; 15'd29155: duty=92; 15'd29156: duty=101; 15'd29157: duty=112; 15'd29158: duty=98; 15'd29159: duty=99;
15'd29160: duty=101; 15'd29161: duty=90; 15'd29162: duty=121; 15'd29163: duty=127; 15'd29164: duty=125; 15'd29165: duty=121; 15'd29166: duty=119; 15'd29167: duty=126;
15'd29168: duty=124; 15'd29169: duty=137; 15'd29170: duty=128; 15'd29171: duty=126; 15'd29172: duty=131; 15'd29173: duty=131; 15'd29174: duty=136; 15'd29175: duty=136;
15'd29176: duty=148; 15'd29177: duty=132; 15'd29178: duty=126; 15'd29179: duty=134; 15'd29180: duty=126; 15'd29181: duty=132; 15'd29182: duty=136; 15'd29183: duty=137;
15'd29184: duty=148; 15'd29185: duty=154; 15'd29186: duty=160; 15'd29187: duty=165; 15'd29188: duty=164; 15'd29189: duty=168; 15'd29190: duty=158; 15'd29191: duty=153;
15'd29192: duty=150; 15'd29193: duty=146; 15'd29194: duty=146; 15'd29195: duty=157; 15'd29196: duty=158; 15'd29197: duty=162; 15'd29198: duty=157; 15'd29199: duty=155;
15'd29200: duty=151; 15'd29201: duty=143; 15'd29202: duty=165; 15'd29203: duty=162; 15'd29204: duty=145; 15'd29205: duty=142; 15'd29206: duty=148; 15'd29207: duty=130;
15'd29208: duty=133; 15'd29209: duty=124; 15'd29210: duty=123; 15'd29211: duty=133; 15'd29212: duty=128; 15'd29213: duty=138; 15'd29214: duty=146; 15'd29215: duty=143;
15'd29216: duty=134; 15'd29217: duty=137; 15'd29218: duty=130; 15'd29219: duty=132; 15'd29220: duty=119; 15'd29221: duty=103; 15'd29222: duty=91; 15'd29223: duty=92;
15'd29224: duty=106; 15'd29225: duty=87; 15'd29226: duty=102; 15'd29227: duty=103; 15'd29228: duty=92; 15'd29229: duty=105; 15'd29230: duty=111; 15'd29231: duty=103;
15'd29232: duty=109; 15'd29233: duty=111; 15'd29234: duty=90; 15'd29235: duty=109; 15'd29236: duty=121; 15'd29237: duty=124; 15'd29238: duty=134; 15'd29239: duty=128;
15'd29240: duty=128; 15'd29241: duty=130; 15'd29242: duty=129; 15'd29243: duty=130; 15'd29244: duty=111; 15'd29245: duty=113; 15'd29246: duty=118; 15'd29247: duty=128;
15'd29248: duty=130; 15'd29249: duty=127; 15'd29250: duty=130; 15'd29251: duty=125; 15'd29252: duty=135; 15'd29253: duty=137; 15'd29254: duty=153; 15'd29255: duty=155;
15'd29256: duty=156; 15'd29257: duty=143; 15'd29258: duty=138; 15'd29259: duty=149; 15'd29260: duty=138; 15'd29261: duty=137; 15'd29262: duty=147; 15'd29263: duty=155;
15'd29264: duty=148; 15'd29265: duty=157; 15'd29266: duty=154; 15'd29267: duty=146; 15'd29268: duty=146; 15'd29269: duty=135; 15'd29270: duty=153; 15'd29271: duty=139;
15'd29272: duty=142; 15'd29273: duty=137; 15'd29274: duty=115; 15'd29275: duty=116; 15'd29276: duty=125; 15'd29277: duty=124; 15'd29278: duty=124; 15'd29279: duty=131;
15'd29280: duty=107; 15'd29281: duty=124; 15'd29282: duty=127; 15'd29283: duty=121; 15'd29284: duty=125; 15'd29285: duty=128; 15'd29286: duty=128; 15'd29287: duty=128;
15'd29288: duty=122; 15'd29289: duty=123; 15'd29290: duty=116; 15'd29291: duty=108; 15'd29292: duty=114; 15'd29293: duty=111; 15'd29294: duty=111; 15'd29295: duty=115;
15'd29296: duty=118; 15'd29297: duty=120; 15'd29298: duty=135; 15'd29299: duty=130; 15'd29300: duty=137; 15'd29301: duty=140; 15'd29302: duty=124; 15'd29303: duty=132;
15'd29304: duty=138; 15'd29305: duty=136; 15'd29306: duty=128; 15'd29307: duty=125; 15'd29308: duty=134; 15'd29309: duty=132; 15'd29310: duty=141; 15'd29311: duty=141;
15'd29312: duty=154; 15'd29313: duty=152; 15'd29314: duty=152; 15'd29315: duty=153; 15'd29316: duty=152; 15'd29317: duty=142; 15'd29318: duty=140; 15'd29319: duty=139;
15'd29320: duty=124; 15'd29321: duty=126; 15'd29322: duty=117; 15'd29323: duty=136; 15'd29324: duty=131; 15'd29325: duty=137; 15'd29326: duty=151; 15'd29327: duty=140;
15'd29328: duty=136; 15'd29329: duty=141; 15'd29330: duty=154; 15'd29331: duty=148; 15'd29332: duty=148; 15'd29333: duty=142; 15'd29334: duty=121; 15'd29335: duty=131;
15'd29336: duty=142; 15'd29337: duty=147; 15'd29338: duty=134; 15'd29339: duty=124; 15'd29340: duty=131; 15'd29341: duty=123; 15'd29342: duty=135; 15'd29343: duty=134;
15'd29344: duty=128; 15'd29345: duty=120; 15'd29346: duty=129; 15'd29347: duty=124; 15'd29348: duty=105; 15'd29349: duty=114; 15'd29350: duty=103; 15'd29351: duty=121;
15'd29352: duty=122; 15'd29353: duty=110; 15'd29354: duty=126; 15'd29355: duty=127; 15'd29356: duty=123; 15'd29357: duty=132; 15'd29358: duty=124; 15'd29359: duty=113;
15'd29360: duty=124; 15'd29361: duty=118; 15'd29362: duty=126; 15'd29363: duty=123; 15'd29364: duty=109; 15'd29365: duty=114; 15'd29366: duty=108; 15'd29367: duty=109;
15'd29368: duty=110; 15'd29369: duty=106; 15'd29370: duty=101; 15'd29371: duty=105; 15'd29372: duty=122; 15'd29373: duty=121; 15'd29374: duty=118; 15'd29375: duty=108;
15'd29376: duty=119; 15'd29377: duty=124; 15'd29378: duty=126; 15'd29379: duty=131; 15'd29380: duty=135; 15'd29381: duty=150; 15'd29382: duty=154; 15'd29383: duty=154;
15'd29384: duty=152; 15'd29385: duty=148; 15'd29386: duty=140; 15'd29387: duty=141; 15'd29388: duty=135; 15'd29389: duty=136; 15'd29390: duty=132; 15'd29391: duty=125;
15'd29392: duty=131; 15'd29393: duty=140; 15'd29394: duty=143; 15'd29395: duty=143; 15'd29396: duty=148; 15'd29397: duty=148; 15'd29398: duty=148; 15'd29399: duty=150;
15'd29400: duty=160; 15'd29401: duty=164; 15'd29402: duty=152; 15'd29403: duty=151; 15'd29404: duty=158; 15'd29405: duty=160; 15'd29406: duty=157; 15'd29407: duty=145;
15'd29408: duty=145; 15'd29409: duty=137; 15'd29410: duty=134; 15'd29411: duty=150; 15'd29412: duty=153; 15'd29413: duty=148; 15'd29414: duty=141; 15'd29415: duty=135;
15'd29416: duty=138; 15'd29417: duty=137; 15'd29418: duty=130; 15'd29419: duty=133; 15'd29420: duty=128; 15'd29421: duty=124; 15'd29422: duty=121; 15'd29423: duty=115;
15'd29424: duty=115; 15'd29425: duty=99; 15'd29426: duty=118; 15'd29427: duty=113; 15'd29428: duty=122; 15'd29429: duty=123; 15'd29430: duty=107; 15'd29431: duty=113;
15'd29432: duty=108; 15'd29433: duty=106; 15'd29434: duty=109; 15'd29435: duty=112; 15'd29436: duty=104; 15'd29437: duty=115; 15'd29438: duty=110; 15'd29439: duty=119;
15'd29440: duty=121; 15'd29441: duty=124; 15'd29442: duty=121; 15'd29443: duty=112; 15'd29444: duty=113; 15'd29445: duty=117; 15'd29446: duty=120; 15'd29447: duty=121;
15'd29448: duty=118; 15'd29449: duty=112; 15'd29450: duty=109; 15'd29451: duty=115; 15'd29452: duty=119; 15'd29453: duty=134; 15'd29454: duty=139; 15'd29455: duty=142;
15'd29456: duty=151; 15'd29457: duty=151; 15'd29458: duty=149; 15'd29459: duty=133; 15'd29460: duty=119; 15'd29461: duty=121; 15'd29462: duty=130; 15'd29463: duty=131;
15'd29464: duty=137; 15'd29465: duty=136; 15'd29466: duty=137; 15'd29467: duty=142; 15'd29468: duty=148; 15'd29469: duty=146; 15'd29470: duty=158; 15'd29471: duty=153;
15'd29472: duty=158; 15'd29473: duty=168; 15'd29474: duty=160; 15'd29475: duty=156; 15'd29476: duty=156; 15'd29477: duty=142; 15'd29478: duty=139; 15'd29479: duty=142;
15'd29480: duty=145; 15'd29481: duty=153; 15'd29482: duty=156; 15'd29483: duty=150; 15'd29484: duty=140; 15'd29485: duty=134; 15'd29486: duty=128; 15'd29487: duty=130;
15'd29488: duty=127; 15'd29489: duty=128; 15'd29490: duty=128; 15'd29491: duty=130; 15'd29492: duty=116; 15'd29493: duty=113; 15'd29494: duty=119; 15'd29495: duty=115;
15'd29496: duty=107; 15'd29497: duty=102; 15'd29498: duty=104; 15'd29499: duty=116; 15'd29500: duty=124; 15'd29501: duty=117; 15'd29502: duty=115; 15'd29503: duty=110;
15'd29504: duty=98; 15'd29505: duty=119; 15'd29506: duty=115; 15'd29507: duty=111; 15'd29508: duty=110; 15'd29509: duty=97; 15'd29510: duty=100; 15'd29511: duty=105;
15'd29512: duty=109; 15'd29513: duty=111; 15'd29514: duty=111; 15'd29515: duty=111; 15'd29516: duty=121; 15'd29517: duty=113; 15'd29518: duty=120; 15'd29519: duty=122;
15'd29520: duty=123; 15'd29521: duty=121; 15'd29522: duty=136; 15'd29523: duty=148; 15'd29524: duty=133; 15'd29525: duty=136; 15'd29526: duty=133; 15'd29527: duty=149;
15'd29528: duty=145; 15'd29529: duty=134; 15'd29530: duty=146; 15'd29531: duty=149; 15'd29532: duty=151; 15'd29533: duty=156; 15'd29534: duty=146; 15'd29535: duty=148;
15'd29536: duty=151; 15'd29537: duty=156; 15'd29538: duty=154; 15'd29539: duty=145; 15'd29540: duty=154; 15'd29541: duty=155; 15'd29542: duty=161; 15'd29543: duty=157;
15'd29544: duty=165; 15'd29545: duty=159; 15'd29546: duty=157; 15'd29547: duty=152; 15'd29548: duty=166; 15'd29549: duty=162; 15'd29550: duty=169; 15'd29551: duty=165;
15'd29552: duty=148; 15'd29553: duty=162; 15'd29554: duty=145; 15'd29555: duty=142; 15'd29556: duty=145; 15'd29557: duty=137; 15'd29558: duty=126; 15'd29559: duty=125;
15'd29560: duty=129; 15'd29561: duty=140; 15'd29562: duty=135; 15'd29563: duty=136; 15'd29564: duty=115; 15'd29565: duty=107; 15'd29566: duty=110; 15'd29567: duty=102;
15'd29568: duty=109; 15'd29569: duty=105; 15'd29570: duty=110; 15'd29571: duty=109; 15'd29572: duty=106; 15'd29573: duty=117; 15'd29574: duty=116; 15'd29575: duty=101;
15'd29576: duty=89; 15'd29577: duty=86; 15'd29578: duty=92; 15'd29579: duty=96; 15'd29580: duty=92; 15'd29581: duty=93; 15'd29582: duty=91; 15'd29583: duty=100;
15'd29584: duty=115; 15'd29585: duty=104; 15'd29586: duty=110; 15'd29587: duty=119; 15'd29588: duty=107; 15'd29589: duty=116; 15'd29590: duty=120; 15'd29591: duty=127;
15'd29592: duty=125; 15'd29593: duty=122; 15'd29594: duty=139; 15'd29595: duty=141; 15'd29596: duty=136; 15'd29597: duty=148; 15'd29598: duty=153; 15'd29599: duty=157;
15'd29600: duty=167; 15'd29601: duty=162; 15'd29602: duty=169; 15'd29603: duty=154; 15'd29604: duty=149; 15'd29605: duty=143; 15'd29606: duty=135; 15'd29607: duty=127;
15'd29608: duty=124; 15'd29609: duty=134; 15'd29610: duty=128; 15'd29611: duty=131; 15'd29612: duty=144; 15'd29613: duty=157; 15'd29614: duty=153; 15'd29615: duty=163;
15'd29616: duty=161; 15'd29617: duty=156; 15'd29618: duty=154; 15'd29619: duty=148; 15'd29620: duty=154; 15'd29621: duty=151; 15'd29622: duty=144; 15'd29623: duty=148;
15'd29624: duty=147; 15'd29625: duty=138; 15'd29626: duty=137; 15'd29627: duty=136; 15'd29628: duty=132; 15'd29629: duty=140; 15'd29630: duty=146; 15'd29631: duty=136;
15'd29632: duty=129; 15'd29633: duty=119; 15'd29634: duty=114; 15'd29635: duty=121; 15'd29636: duty=113; 15'd29637: duty=115; 15'd29638: duty=108; 15'd29639: duty=115;
15'd29640: duty=116; 15'd29641: duty=112; 15'd29642: duty=123; 15'd29643: duty=115; 15'd29644: duty=113; 15'd29645: duty=107; 15'd29646: duty=118; 15'd29647: duty=120;
15'd29648: duty=125; 15'd29649: duty=90; 15'd29650: duty=87; 15'd29651: duty=105; 15'd29652: duty=95; 15'd29653: duty=102; 15'd29654: duty=109; 15'd29655: duty=113;
15'd29656: duty=112; 15'd29657: duty=121; 15'd29658: duty=109; 15'd29659: duty=108; 15'd29660: duty=104; 15'd29661: duty=88; 15'd29662: duty=93; 15'd29663: duty=113;
15'd29664: duty=121; 15'd29665: duty=125; 15'd29666: duty=120; 15'd29667: duty=137; 15'd29668: duty=152; 15'd29669: duty=142; 15'd29670: duty=133; 15'd29671: duty=142;
15'd29672: duty=160; 15'd29673: duty=154; 15'd29674: duty=153; 15'd29675: duty=160; 15'd29676: duty=150; 15'd29677: duty=152; 15'd29678: duty=158; 15'd29679: duty=154;
15'd29680: duty=170; 15'd29681: duty=172; 15'd29682: duty=169; 15'd29683: duty=176; 15'd29684: duty=173; 15'd29685: duty=176; 15'd29686: duty=170; 15'd29687: duty=166;
15'd29688: duty=159; 15'd29689: duty=153; 15'd29690: duty=165; 15'd29691: duty=168; 15'd29692: duty=162; 15'd29693: duty=156; 15'd29694: duty=155; 15'd29695: duty=157;
15'd29696: duty=159; 15'd29697: duty=153; 15'd29698: duty=148; 15'd29699: duty=142; 15'd29700: duty=143; 15'd29701: duty=133; 15'd29702: duty=134; 15'd29703: duty=138;
15'd29704: duty=132; 15'd29705: duty=121; 15'd29706: duty=120; 15'd29707: duty=115; 15'd29708: duty=117; 15'd29709: duty=112; 15'd29710: duty=94; 15'd29711: duty=97;
15'd29712: duty=93; 15'd29713: duty=95; 15'd29714: duty=93; 15'd29715: duty=99; 15'd29716: duty=100; 15'd29717: duty=101; 15'd29718: duty=108; 15'd29719: duty=95;
15'd29720: duty=97; 15'd29721: duty=102; 15'd29722: duty=85; 15'd29723: duty=95; 15'd29724: duty=87; 15'd29725: duty=89; 15'd29726: duty=99; 15'd29727: duty=84;
15'd29728: duty=93; 15'd29729: duty=101; 15'd29730: duty=106; 15'd29731: duty=110; 15'd29732: duty=106; 15'd29733: duty=99; 15'd29734: duty=101; 15'd29735: duty=121;
15'd29736: duty=120; 15'd29737: duty=115; 15'd29738: duty=121; 15'd29739: duty=128; 15'd29740: duty=143; 15'd29741: duty=143; 15'd29742: duty=138; 15'd29743: duty=138;
15'd29744: duty=144; 15'd29745: duty=160; 15'd29746: duty=153; 15'd29747: duty=151; 15'd29748: duty=146; 15'd29749: duty=140; 15'd29750: duty=138; 15'd29751: duty=143;
15'd29752: duty=136; 15'd29753: duty=143; 15'd29754: duty=152; 15'd29755: duty=151; 15'd29756: duty=169; 15'd29757: duty=177; 15'd29758: duty=184; 15'd29759: duty=180;
15'd29760: duty=172; 15'd29761: duty=161; 15'd29762: duty=165; 15'd29763: duty=161; 15'd29764: duty=161; 15'd29765: duty=158; 15'd29766: duty=161; 15'd29767: duty=166;
15'd29768: duty=166; 15'd29769: duty=170; 15'd29770: duty=160; 15'd29771: duty=164; 15'd29772: duty=171; 15'd29773: duty=157; 15'd29774: duty=161; 15'd29775: duty=152;
15'd29776: duty=142; 15'd29777: duty=143; 15'd29778: duty=140; 15'd29779: duty=135; 15'd29780: duty=113; 15'd29781: duty=110; 15'd29782: duty=104; 15'd29783: duty=110;
15'd29784: duty=118; 15'd29785: duty=140; 15'd29786: duty=120; 15'd29787: duty=118; 15'd29788: duty=112; 15'd29789: duty=90; 15'd29790: duty=101; 15'd29791: duty=90;
15'd29792: duty=97; 15'd29793: duty=94; 15'd29794: duty=89; 15'd29795: duty=82; 15'd29796: duty=78; 15'd29797: duty=91; 15'd29798: duty=83; 15'd29799: duty=84;
15'd29800: duty=97; 15'd29801: duty=102; 15'd29802: duty=114; 15'd29803: duty=115; 15'd29804: duty=93; 15'd29805: duty=97; 15'd29806: duty=105; 15'd29807: duty=100;
15'd29808: duty=100; 15'd29809: duty=102; 15'd29810: duty=101; 15'd29811: duty=101; 15'd29812: duty=115; 15'd29813: duty=123; 15'd29814: duty=128; 15'd29815: duty=128;
15'd29816: duty=139; 15'd29817: duty=124; 15'd29818: duty=127; 15'd29819: duty=141; 15'd29820: duty=144; 15'd29821: duty=149; 15'd29822: duty=136; 15'd29823: duty=143;
15'd29824: duty=150; 15'd29825: duty=151; 15'd29826: duty=149; 15'd29827: duty=160; 15'd29828: duty=165; 15'd29829: duty=168; 15'd29830: duty=159; 15'd29831: duty=172;
15'd29832: duty=174; 15'd29833: duty=165; 15'd29834: duty=171; 15'd29835: duty=169; 15'd29836: duty=176; 15'd29837: duty=185; 15'd29838: duty=176; 15'd29839: duty=173;
15'd29840: duty=172; 15'd29841: duty=156; 15'd29842: duty=156; 15'd29843: duty=167; 15'd29844: duty=151; 15'd29845: duty=141; 15'd29846: duty=147; 15'd29847: duty=136;
15'd29848: duty=136; 15'd29849: duty=121; 15'd29850: duty=129; 15'd29851: duty=127; 15'd29852: duty=108; 15'd29853: duty=120; 15'd29854: duty=114; 15'd29855: duty=112;
15'd29856: duty=121; 15'd29857: duty=107; 15'd29858: duty=113; 15'd29859: duty=112; 15'd29860: duty=111; 15'd29861: duty=119; 15'd29862: duty=106; 15'd29863: duty=97;
15'd29864: duty=95; 15'd29865: duty=102; 15'd29866: duty=110; 15'd29867: duty=116; 15'd29868: duty=105; 15'd29869: duty=106; 15'd29870: duty=108; 15'd29871: duty=107;
15'd29872: duty=99; 15'd29873: duty=103; 15'd29874: duty=96; 15'd29875: duty=99; 15'd29876: duty=107; 15'd29877: duty=114; 15'd29878: duty=125; 15'd29879: duty=130;
15'd29880: duty=132; 15'd29881: duty=128; 15'd29882: duty=133; 15'd29883: duty=140; 15'd29884: duty=145; 15'd29885: duty=148; 15'd29886: duty=146; 15'd29887: duty=142;
15'd29888: duty=154; 15'd29889: duty=157; 15'd29890: duty=160; 15'd29891: duty=139; 15'd29892: duty=128; 15'd29893: duty=133; 15'd29894: duty=140; 15'd29895: duty=136;
15'd29896: duty=143; 15'd29897: duty=151; 15'd29898: duty=145; 15'd29899: duty=146; 15'd29900: duty=142; 15'd29901: duty=146; 15'd29902: duty=153; 15'd29903: duty=159;
15'd29904: duty=160; 15'd29905: duty=168; 15'd29906: duty=162; 15'd29907: duty=160; 15'd29908: duty=151; 15'd29909: duty=143; 15'd29910: duty=145; 15'd29911: duty=140;
15'd29912: duty=145; 15'd29913: duty=147; 15'd29914: duty=153; 15'd29915: duty=140; 15'd29916: duty=131; 15'd29917: duty=128; 15'd29918: duty=134; 15'd29919: duty=140;
15'd29920: duty=117; 15'd29921: duty=109; 15'd29922: duty=108; 15'd29923: duty=111; 15'd29924: duty=119; 15'd29925: duty=117; 15'd29926: duty=116; 15'd29927: duty=123;
15'd29928: duty=113; 15'd29929: duty=110; 15'd29930: duty=131; 15'd29931: duty=123; 15'd29932: duty=116; 15'd29933: duty=127; 15'd29934: duty=98; 15'd29935: duty=89;
15'd29936: duty=91; 15'd29937: duty=87; 15'd29938: duty=77; 15'd29939: duty=94; 15'd29940: duty=111; 15'd29941: duty=102; 15'd29942: duty=97; 15'd29943: duty=94;
15'd29944: duty=103; 15'd29945: duty=126; 15'd29946: duty=123; 15'd29947: duty=100; 15'd29948: duty=99; 15'd29949: duty=106; 15'd29950: duty=126; 15'd29951: duty=143;
15'd29952: duty=139; 15'd29953: duty=141; 15'd29954: duty=143; 15'd29955: duty=123; 15'd29956: duty=140; 15'd29957: duty=124; 15'd29958: duty=125; 15'd29959: duty=131;
15'd29960: duty=117; 15'd29961: duty=133; 15'd29962: duty=128; 15'd29963: duty=136; 15'd29964: duty=139; 15'd29965: duty=128; 15'd29966: duty=146; 15'd29967: duty=145;
15'd29968: duty=154; 15'd29969: duty=165; 15'd29970: duty=166; 15'd29971: duty=169; 15'd29972: duty=161; 15'd29973: duty=158; 15'd29974: duty=166; 15'd29975: duty=159;
15'd29976: duty=163; 15'd29977: duty=165; 15'd29978: duty=154; 15'd29979: duty=160; 15'd29980: duty=151; 15'd29981: duty=152; 15'd29982: duty=158; 15'd29983: duty=146;
15'd29984: duty=152; 15'd29985: duty=166; 15'd29986: duty=155; 15'd29987: duty=162; 15'd29988: duty=159; 15'd29989: duty=166; 15'd29990: duty=141; 15'd29991: duty=133;
15'd29992: duty=112; 15'd29993: duty=113; 15'd29994: duty=139; 15'd29995: duty=132; 15'd29996: duty=124; 15'd29997: duty=135; 15'd29998: duty=131; 15'd29999: duty=129;
15'd30000: duty=137; 15'd30001: duty=120; 15'd30002: duty=112; 15'd30003: duty=113; 15'd30004: duty=123; 15'd30005: duty=113; 15'd30006: duty=118; 15'd30007: duty=99;
15'd30008: duty=91; 15'd30009: duty=96; 15'd30010: duty=99; 15'd30011: duty=112; 15'd30012: duty=112; 15'd30013: duty=101; 15'd30014: duty=99; 15'd30015: duty=104;
15'd30016: duty=114; 15'd30017: duty=129; 15'd30018: duty=128; 15'd30019: duty=98; 15'd30020: duty=102; 15'd30021: duty=95; 15'd30022: duty=118; 15'd30023: duty=126;
15'd30024: duty=111; 15'd30025: duty=118; 15'd30026: duty=117; 15'd30027: duty=133; 15'd30028: duty=146; 15'd30029: duty=142; 15'd30030: duty=127; 15'd30031: duty=126;
15'd30032: duty=124; 15'd30033: duty=122; 15'd30034: duty=127; 15'd30035: duty=133; 15'd30036: duty=127; 15'd30037: duty=121; 15'd30038: duty=113; 15'd30039: duty=124;
15'd30040: duty=127; 15'd30041: duty=138; 15'd30042: duty=124; 15'd30043: duty=139; 15'd30044: duty=157; 15'd30045: duty=156; 15'd30046: duty=160; 15'd30047: duty=140;
15'd30048: duty=145; 15'd30049: duty=148; 15'd30050: duty=151; 15'd30051: duty=149; 15'd30052: duty=151; 15'd30053: duty=162; 15'd30054: duty=167; 15'd30055: duty=172;
15'd30056: duty=170; 15'd30057: duty=168; 15'd30058: duty=156; 15'd30059: duty=150; 15'd30060: duty=137; 15'd30061: duty=141; 15'd30062: duty=135; 15'd30063: duty=129;
15'd30064: duty=137; 15'd30065: duty=135; 15'd30066: duty=148; 15'd30067: duty=145; 15'd30068: duty=136; 15'd30069: duty=120; 15'd30070: duty=113; 15'd30071: duty=119;
15'd30072: duty=124; 15'd30073: duty=119; 15'd30074: duty=124; 15'd30075: duty=117; 15'd30076: duty=109; 15'd30077: duty=106; 15'd30078: duty=107; 15'd30079: duty=102;
15'd30080: duty=89; 15'd30081: duty=99; 15'd30082: duty=116; 15'd30083: duty=113; 15'd30084: duty=104; 15'd30085: duty=96; 15'd30086: duty=98; 15'd30087: duty=94;
15'd30088: duty=99; 15'd30089: duty=102; 15'd30090: duty=95; 15'd30091: duty=102; 15'd30092: duty=106; 15'd30093: duty=112; 15'd30094: duty=110; 15'd30095: duty=105;
15'd30096: duty=106; 15'd30097: duty=113; 15'd30098: duty=118; 15'd30099: duty=127; 15'd30100: duty=133; 15'd30101: duty=139; 15'd30102: duty=129; 15'd30103: duty=127;
15'd30104: duty=123; 15'd30105: duty=119; 15'd30106: duty=138; 15'd30107: duty=146; 15'd30108: duty=141; 15'd30109: duty=148; 15'd30110: duty=141; 15'd30111: duty=143;
15'd30112: duty=163; 15'd30113: duty=160; 15'd30114: duty=163; 15'd30115: duty=169; 15'd30116: duty=176; 15'd30117: duty=177; 15'd30118: duty=176; 15'd30119: duty=177;
15'd30120: duty=178; 15'd30121: duty=187; 15'd30122: duty=185; 15'd30123: duty=178; 15'd30124: duty=182; 15'd30125: duty=194; 15'd30126: duty=181; 15'd30127: duty=172;
15'd30128: duty=166; 15'd30129: duty=158; 15'd30130: duty=164; 15'd30131: duty=146; 15'd30132: duty=147; 15'd30133: duty=141; 15'd30134: duty=141; 15'd30135: duty=140;
15'd30136: duty=145; 15'd30137: duty=141; 15'd30138: duty=137; 15'd30139: duty=125; 15'd30140: duty=101; 15'd30141: duty=117; 15'd30142: duty=96; 15'd30143: duty=101;
15'd30144: duty=112; 15'd30145: duty=99; 15'd30146: duty=108; 15'd30147: duty=104; 15'd30148: duty=98; 15'd30149: duty=98; 15'd30150: duty=92; 15'd30151: duty=90;
15'd30152: duty=87; 15'd30153: duty=87; 15'd30154: duty=97; 15'd30155: duty=101; 15'd30156: duty=82; 15'd30157: duty=84; 15'd30158: duty=84; 15'd30159: duty=86;
15'd30160: duty=100; 15'd30161: duty=107; 15'd30162: duty=107; 15'd30163: duty=101; 15'd30164: duty=104; 15'd30165: duty=112; 15'd30166: duty=115; 15'd30167: duty=121;
15'd30168: duty=113; 15'd30169: duty=107; 15'd30170: duty=124; 15'd30171: duty=134; 15'd30172: duty=129; 15'd30173: duty=121; 15'd30174: duty=131; 15'd30175: duty=129;
15'd30176: duty=140; 15'd30177: duty=135; 15'd30178: duty=122; 15'd30179: duty=124; 15'd30180: duty=121; 15'd30181: duty=126; 15'd30182: duty=139; 15'd30183: duty=139;
15'd30184: duty=154; 15'd30185: duty=159; 15'd30186: duty=149; 15'd30187: duty=160; 15'd30188: duty=168; 15'd30189: duty=168; 15'd30190: duty=172; 15'd30191: duty=154;
15'd30192: duty=150; 15'd30193: duty=163; 15'd30194: duty=166; 15'd30195: duty=160; 15'd30196: duty=171; 15'd30197: duty=168; 15'd30198: duty=137; 15'd30199: duty=141;
15'd30200: duty=140; 15'd30201: duty=154; 15'd30202: duty=171; 15'd30203: duty=162; 15'd30204: duty=151; 15'd30205: duty=141; 15'd30206: duty=131; 15'd30207: duty=145;
15'd30208: duty=128; 15'd30209: duty=121; 15'd30210: duty=133; 15'd30211: duty=133; 15'd30212: duty=132; 15'd30213: duty=122; 15'd30214: duty=121; 15'd30215: duty=135;
15'd30216: duty=131; 15'd30217: duty=120; 15'd30218: duty=122; 15'd30219: duty=109; 15'd30220: duty=115; 15'd30221: duty=112; 15'd30222: duty=117; 15'd30223: duty=119;
15'd30224: duty=91; 15'd30225: duty=97; 15'd30226: duty=101; 15'd30227: duty=104; 15'd30228: duty=123; 15'd30229: duty=112; 15'd30230: duty=107; 15'd30231: duty=114;
15'd30232: duty=111; 15'd30233: duty=115; 15'd30234: duty=122; 15'd30235: duty=115; 15'd30236: duty=122; 15'd30237: duty=120; 15'd30238: duty=129; 15'd30239: duty=130;
15'd30240: duty=134; 15'd30241: duty=141; 15'd30242: duty=129; 15'd30243: duty=125; 15'd30244: duty=128; 15'd30245: duty=132; 15'd30246: duty=131; 15'd30247: duty=129;
15'd30248: duty=131; 15'd30249: duty=141; 15'd30250: duty=140; 15'd30251: duty=144; 15'd30252: duty=137; 15'd30253: duty=147; 15'd30254: duty=160; 15'd30255: duty=161;
15'd30256: duty=151; 15'd30257: duty=142; 15'd30258: duty=142; 15'd30259: duty=147; 15'd30260: duty=143; 15'd30261: duty=154; 15'd30262: duty=151; 15'd30263: duty=147;
15'd30264: duty=146; 15'd30265: duty=139; 15'd30266: duty=149; 15'd30267: duty=154; 15'd30268: duty=158; 15'd30269: duty=153; 15'd30270: duty=145; 15'd30271: duty=145;
15'd30272: duty=145; 15'd30273: duty=133; 15'd30274: duty=136; 15'd30275: duty=133; 15'd30276: duty=132; 15'd30277: duty=122; 15'd30278: duty=121; 15'd30279: duty=128;
15'd30280: duty=119; 15'd30281: duty=114; 15'd30282: duty=112; 15'd30283: duty=125; 15'd30284: duty=127; 15'd30285: duty=107; 15'd30286: duty=98; 15'd30287: duty=105;
15'd30288: duty=106; 15'd30289: duty=100; 15'd30290: duty=108; 15'd30291: duty=96; 15'd30292: duty=107; 15'd30293: duty=115; 15'd30294: duty=109; 15'd30295: duty=107;
15'd30296: duty=97; 15'd30297: duty=101; 15'd30298: duty=98; 15'd30299: duty=105; 15'd30300: duty=106; 15'd30301: duty=110; 15'd30302: duty=108; 15'd30303: duty=107;
15'd30304: duty=114; 15'd30305: duty=121; 15'd30306: duty=114; 15'd30307: duty=110; 15'd30308: duty=108; 15'd30309: duty=126; 15'd30310: duty=138; 15'd30311: duty=141;
15'd30312: duty=140; 15'd30313: duty=127; 15'd30314: duty=141; 15'd30315: duty=128; 15'd30316: duty=132; 15'd30317: duty=146; 15'd30318: duty=136; 15'd30319: duty=160;
15'd30320: duty=161; 15'd30321: duty=157; 15'd30322: duty=150; 15'd30323: duty=159; 15'd30324: duty=153; 15'd30325: duty=146; 15'd30326: duty=138; 15'd30327: duty=138;
15'd30328: duty=148; 15'd30329: duty=149; 15'd30330: duty=175; 15'd30331: duty=162; 15'd30332: duty=147; 15'd30333: duty=157; 15'd30334: duty=173; 15'd30335: duty=174;
15'd30336: duty=184; 15'd30337: duty=177; 15'd30338: duty=159; 15'd30339: duty=154; 15'd30340: duty=159; 15'd30341: duty=156; 15'd30342: duty=156; 15'd30343: duty=144;
15'd30344: duty=144; 15'd30345: duty=140; 15'd30346: duty=134; 15'd30347: duty=150; 15'd30348: duty=145; 15'd30349: duty=127; 15'd30350: duty=136; 15'd30351: duty=139;
15'd30352: duty=141; 15'd30353: duty=150; 15'd30354: duty=121; 15'd30355: duty=116; 15'd30356: duty=112; 15'd30357: duty=106; 15'd30358: duty=113; 15'd30359: duty=116;
15'd30360: duty=131; 15'd30361: duty=113; 15'd30362: duty=98; 15'd30363: duty=94; 15'd30364: duty=96; 15'd30365: duty=101; 15'd30366: duty=99; 15'd30367: duty=107;
15'd30368: duty=96; 15'd30369: duty=102; 15'd30370: duty=92; 15'd30371: duty=96; 15'd30372: duty=101; 15'd30373: duty=111; 15'd30374: duty=99; 15'd30375: duty=83;
15'd30376: duty=86; 15'd30377: duty=104; 15'd30378: duty=124; 15'd30379: duty=116; 15'd30380: duty=110; 15'd30381: duty=117; 15'd30382: duty=128; 15'd30383: duty=124;
15'd30384: duty=111; 15'd30385: duty=107; 15'd30386: duty=107; 15'd30387: duty=106; 15'd30388: duty=112; 15'd30389: duty=104; 15'd30390: duty=108; 15'd30391: duty=118;
15'd30392: duty=135; 15'd30393: duty=142; 15'd30394: duty=137; 15'd30395: duty=135; 15'd30396: duty=139; 15'd30397: duty=144; 15'd30398: duty=148; 15'd30399: duty=148;
15'd30400: duty=159; 15'd30401: duty=149; 15'd30402: duty=143; 15'd30403: duty=155; 15'd30404: duty=165; 15'd30405: duty=161; 15'd30406: duty=157; 15'd30407: duty=162;
15'd30408: duty=168; 15'd30409: duty=179; 15'd30410: duty=168; 15'd30411: duty=167; 15'd30412: duty=157; 15'd30413: duty=148; 15'd30414: duty=145; 15'd30415: duty=147;
15'd30416: duty=149; 15'd30417: duty=141; 15'd30418: duty=142; 15'd30419: duty=142; 15'd30420: duty=143; 15'd30421: duty=139; 15'd30422: duty=164; 15'd30423: duty=136;
15'd30424: duty=132; 15'd30425: duty=154; 15'd30426: duty=123; 15'd30427: duty=136; 15'd30428: duty=128; 15'd30429: duty=125; 15'd30430: duty=129; 15'd30431: duty=122;
15'd30432: duty=127; 15'd30433: duty=125; 15'd30434: duty=128; 15'd30435: duty=124; 15'd30436: duty=112; 15'd30437: duty=101; 15'd30438: duty=95; 15'd30439: duty=110;
15'd30440: duty=108; 15'd30441: duty=113; 15'd30442: duty=114; 15'd30443: duty=127; 15'd30444: duty=127; 15'd30445: duty=114; 15'd30446: duty=124; 15'd30447: duty=126;
15'd30448: duty=124; 15'd30449: duty=121; 15'd30450: duty=132; 15'd30451: duty=144; 15'd30452: duty=134; 15'd30453: duty=127; 15'd30454: duty=126; 15'd30455: duty=130;
15'd30456: duty=142; 15'd30457: duty=136; 15'd30458: duty=137; 15'd30459: duty=147; 15'd30460: duty=148; 15'd30461: duty=143; 15'd30462: duty=130; 15'd30463: duty=120;
15'd30464: duty=124; 15'd30465: duty=121; 15'd30466: duty=129; 15'd30467: duty=128; 15'd30468: duty=131; 15'd30469: duty=138; 15'd30470: duty=142; 15'd30471: duty=151;
15'd30472: duty=163; 15'd30473: duty=161; 15'd30474: duty=157; 15'd30475: duty=159; 15'd30476: duty=154; 15'd30477: duty=148; 15'd30478: duty=151; 15'd30479: duty=136;
15'd30480: duty=131; 15'd30481: duty=127; 15'd30482: duty=119; 15'd30483: duty=130; 15'd30484: duty=128; 15'd30485: duty=135; 15'd30486: duty=128; 15'd30487: duty=104;
15'd30488: duty=102; 15'd30489: duty=116; 15'd30490: duty=125; 15'd30491: duty=128; 15'd30492: duty=113; 15'd30493: duty=98; 15'd30494: duty=94; 15'd30495: duty=99;
15'd30496: duty=92; 15'd30497: duty=88; 15'd30498: duty=94; 15'd30499: duty=94; 15'd30500: duty=95; 15'd30501: duty=101; 15'd30502: duty=96; 15'd30503: duty=104;
15'd30504: duty=113; 15'd30505: duty=109; 15'd30506: duty=96; 15'd30507: duty=104; 15'd30508: duty=114; 15'd30509: duty=103; 15'd30510: duty=109; 15'd30511: duty=126;
15'd30512: duty=119; 15'd30513: duty=128; 15'd30514: duty=123; 15'd30515: duty=120; 15'd30516: duty=127; 15'd30517: duty=130; 15'd30518: duty=124; 15'd30519: duty=110;
15'd30520: duty=138; 15'd30521: duty=143; 15'd30522: duty=143; 15'd30523: duty=144; 15'd30524: duty=149; 15'd30525: duty=151; 15'd30526: duty=145; 15'd30527: duty=156;
15'd30528: duty=150; 15'd30529: duty=154; 15'd30530: duty=169; 15'd30531: duty=156; 15'd30532: duty=177; 15'd30533: duty=174; 15'd30534: duty=166; 15'd30535: duty=168;
15'd30536: duty=175; 15'd30537: duty=184; 15'd30538: duty=185; 15'd30539: duty=182; 15'd30540: duty=174; 15'd30541: duty=166; 15'd30542: duty=168; 15'd30543: duty=176;
15'd30544: duty=166; 15'd30545: duty=166; 15'd30546: duty=165; 15'd30547: duty=170; 15'd30548: duty=175; 15'd30549: duty=165; 15'd30550: duty=164; 15'd30551: duty=159;
15'd30552: duty=140; 15'd30553: duty=137; 15'd30554: duty=138; 15'd30555: duty=138; 15'd30556: duty=122; 15'd30557: duty=128; 15'd30558: duty=126; 15'd30559: duty=129;
15'd30560: duty=119; 15'd30561: duty=111; 15'd30562: duty=103; 15'd30563: duty=94; 15'd30564: duty=100; 15'd30565: duty=102; 15'd30566: duty=109; 15'd30567: duty=99;
15'd30568: duty=81; 15'd30569: duty=82; 15'd30570: duty=86; 15'd30571: duty=91; 15'd30572: duty=93; 15'd30573: duty=85; 15'd30574: duty=86; 15'd30575: duty=78;
15'd30576: duty=89; 15'd30577: duty=88; 15'd30578: duty=81; 15'd30579: duty=79; 15'd30580: duty=71; 15'd30581: duty=87; 15'd30582: duty=104; 15'd30583: duty=106;
15'd30584: duty=99; 15'd30585: duty=81; 15'd30586: duty=87; 15'd30587: duty=100; 15'd30588: duty=102; 15'd30589: duty=108; 15'd30590: duty=113; 15'd30591: duty=126;
15'd30592: duty=124; 15'd30593: duty=131; 15'd30594: duty=137; 15'd30595: duty=130; 15'd30596: duty=149; 15'd30597: duty=147; 15'd30598: duty=132; 15'd30599: duty=130;
15'd30600: duty=148; 15'd30601: duty=151; 15'd30602: duty=155; 15'd30603: duty=168; 15'd30604: duty=166; 15'd30605: duty=158; 15'd30606: duty=154; 15'd30607: duty=156;
15'd30608: duty=165; 15'd30609: duty=164; 15'd30610: duty=162; 15'd30611: duty=155; 15'd30612: duty=164; 15'd30613: duty=187; 15'd30614: duty=177; 15'd30615: duty=179;
15'd30616: duty=176; 15'd30617: duty=171; 15'd30618: duty=159; 15'd30619: duty=163; 15'd30620: duty=185; 15'd30621: duty=179; 15'd30622: duty=176; 15'd30623: duty=188;
15'd30624: duty=157; 15'd30625: duty=168; 15'd30626: duty=174; 15'd30627: duty=154; 15'd30628: duty=143; 15'd30629: duty=127; 15'd30630: duty=145; 15'd30631: duty=148;
15'd30632: duty=138; 15'd30633: duty=122; 15'd30634: duty=126; 15'd30635: duty=111; 15'd30636: duty=101; 15'd30637: duty=121; 15'd30638: duty=124; 15'd30639: duty=108;
15'd30640: duty=111; 15'd30641: duty=114; 15'd30642: duty=101; 15'd30643: duty=117; 15'd30644: duty=112; 15'd30645: duty=92; 15'd30646: duty=81; 15'd30647: duty=86;
15'd30648: duty=101; 15'd30649: duty=103; 15'd30650: duty=96; 15'd30651: duty=82; 15'd30652: duty=94; 15'd30653: duty=116; 15'd30654: duty=103; 15'd30655: duty=85;
15'd30656: duty=95; 15'd30657: duty=92; 15'd30658: duty=91; 15'd30659: duty=85; 15'd30660: duty=91; 15'd30661: duty=107; 15'd30662: duty=114; 15'd30663: duty=119;
15'd30664: duty=120; 15'd30665: duty=124; 15'd30666: duty=127; 15'd30667: duty=116; 15'd30668: duty=109; 15'd30669: duty=124; 15'd30670: duty=121; 15'd30671: duty=116;
15'd30672: duty=112; 15'd30673: duty=108; 15'd30674: duty=127; 15'd30675: duty=133; 15'd30676: duty=136; 15'd30677: duty=138; 15'd30678: duty=142; 15'd30679: duty=155;
15'd30680: duty=142; 15'd30681: duty=150; 15'd30682: duty=154; 15'd30683: duty=151; 15'd30684: duty=156; 15'd30685: duty=153; 15'd30686: duty=159; 15'd30687: duty=178;
15'd30688: duty=181; 15'd30689: duty=178; 15'd30690: duty=177; 15'd30691: duty=168; 15'd30692: duty=178; 15'd30693: duty=183; 15'd30694: duty=163; 15'd30695: duty=154;
15'd30696: duty=158; 15'd30697: duty=151; 15'd30698: duty=160; 15'd30699: duty=150; 15'd30700: duty=159; 15'd30701: duty=160; 15'd30702: duty=131; 15'd30703: duty=116;
15'd30704: duty=129; 15'd30705: duty=146; 15'd30706: duty=134; 15'd30707: duty=122; 15'd30708: duty=108; 15'd30709: duty=118; 15'd30710: duty=129; 15'd30711: duty=108;
15'd30712: duty=109; 15'd30713: duty=126; 15'd30714: duty=122; 15'd30715: duty=125; 15'd30716: duty=127; 15'd30717: duty=124; 15'd30718: duty=120; 15'd30719: duty=115;
15'd30720: duty=119; 15'd30721: duty=124; 15'd30722: duty=125; 15'd30723: duty=118; 15'd30724: duty=108; 15'd30725: duty=103; 15'd30726: duty=104; 15'd30727: duty=109;
15'd30728: duty=110; 15'd30729: duty=108; 15'd30730: duty=109; 15'd30731: duty=107; 15'd30732: duty=111; 15'd30733: duty=115; 15'd30734: duty=118; 15'd30735: duty=127;
15'd30736: duty=122; 15'd30737: duty=136; 15'd30738: duty=150; 15'd30739: duty=148; 15'd30740: duty=141; 15'd30741: duty=139; 15'd30742: duty=136; 15'd30743: duty=129;
15'd30744: duty=126; 15'd30745: duty=141; 15'd30746: duty=131; 15'd30747: duty=130; 15'd30748: duty=118; 15'd30749: duty=109; 15'd30750: duty=139; 15'd30751: duty=148;
15'd30752: duty=146; 15'd30753: duty=130; 15'd30754: duty=150; 15'd30755: duty=161; 15'd30756: duty=177; 15'd30757: duty=167; 15'd30758: duty=141; 15'd30759: duty=136;
15'd30760: duty=128; 15'd30761: duty=130; 15'd30762: duty=154; 15'd30763: duty=153; 15'd30764: duty=139; 15'd30765: duty=118; 15'd30766: duty=124; 15'd30767: duty=142;
15'd30768: duty=138; 15'd30769: duty=136; 15'd30770: duty=121; 15'd30771: duty=127; 15'd30772: duty=133; 15'd30773: duty=137; 15'd30774: duty=132; 15'd30775: duty=121;
15'd30776: duty=105; 15'd30777: duty=97; 15'd30778: duty=129; 15'd30779: duty=148; 15'd30780: duty=135; 15'd30781: duty=112; 15'd30782: duty=109; 15'd30783: duty=131;
15'd30784: duty=129; 15'd30785: duty=133; 15'd30786: duty=108; 15'd30787: duty=93; 15'd30788: duty=97; 15'd30789: duty=87; 15'd30790: duty=106; 15'd30791: duty=115;
15'd30792: duty=129; 15'd30793: duty=122; 15'd30794: duty=102; 15'd30795: duty=113; 15'd30796: duty=118; 15'd30797: duty=138; 15'd30798: duty=130; 15'd30799: duty=112;
15'd30800: duty=109; 15'd30801: duty=98; 15'd30802: duty=100; 15'd30803: duty=123; 15'd30804: duty=121; 15'd30805: duty=109; 15'd30806: duty=116; 15'd30807: duty=133;
15'd30808: duty=153; 15'd30809: duty=146; 15'd30810: duty=140; 15'd30811: duty=139; 15'd30812: duty=140; 15'd30813: duty=138; 15'd30814: duty=140; 15'd30815: duty=151;
15'd30816: duty=160; 15'd30817: duty=156; 15'd30818: duty=156; 15'd30819: duty=162; 15'd30820: duty=174; 15'd30821: duty=166; 15'd30822: duty=170; 15'd30823: duty=160;
15'd30824: duty=160; 15'd30825: duty=157; 15'd30826: duty=160; 15'd30827: duty=168; 15'd30828: duty=162; 15'd30829: duty=180; 15'd30830: duty=176; 15'd30831: duty=168;
15'd30832: duty=185; 15'd30833: duty=175; 15'd30834: duty=161; 15'd30835: duty=149; 15'd30836: duty=156; 15'd30837: duty=167; 15'd30838: duty=158; 15'd30839: duty=156;
15'd30840: duty=139; 15'd30841: duty=154; 15'd30842: duty=150; 15'd30843: duty=129; 15'd30844: duty=110; 15'd30845: duty=113; 15'd30846: duty=111; 15'd30847: duty=112;
15'd30848: duty=107; 15'd30849: duty=99; 15'd30850: duty=119; 15'd30851: duty=113; 15'd30852: duty=87; 15'd30853: duty=89; 15'd30854: duty=84; 15'd30855: duty=81;
15'd30856: duty=101; 15'd30857: duty=101; 15'd30858: duty=98; 15'd30859: duty=85; 15'd30860: duty=81; 15'd30861: duty=81; 15'd30862: duty=73; 15'd30863: duty=84;
15'd30864: duty=99; 15'd30865: duty=102; 15'd30866: duty=96; 15'd30867: duty=94; 15'd30868: duty=96; 15'd30869: duty=93; 15'd30870: duty=102; 15'd30871: duty=97;
15'd30872: duty=111; 15'd30873: duty=110; 15'd30874: duty=113; 15'd30875: duty=119; 15'd30876: duty=114; 15'd30877: duty=128; 15'd30878: duty=127; 15'd30879: duty=138;
15'd30880: duty=139; 15'd30881: duty=129; 15'd30882: duty=138; 15'd30883: duty=155; 15'd30884: duty=147; 15'd30885: duty=138; 15'd30886: duty=136; 15'd30887: duty=135;
15'd30888: duty=131; 15'd30889: duty=133; 15'd30890: duty=142; 15'd30891: duty=149; 15'd30892: duty=146; 15'd30893: duty=154; 15'd30894: duty=161; 15'd30895: duty=161;
15'd30896: duty=162; 15'd30897: duty=160; 15'd30898: duty=166; 15'd30899: duty=158; 15'd30900: duty=164; 15'd30901: duty=169; 15'd30902: duty=164; 15'd30903: duty=160;
15'd30904: duty=170; 15'd30905: duty=179; 15'd30906: duty=181; 15'd30907: duty=180; 15'd30908: duty=175; 15'd30909: duty=180; 15'd30910: duty=172; 15'd30911: duty=178;
15'd30912: duty=164; 15'd30913: duty=147; 15'd30914: duty=140; 15'd30915: duty=141; 15'd30916: duty=127; 15'd30917: duty=117; 15'd30918: duty=122; 15'd30919: duty=109;
15'd30920: duty=105; 15'd30921: duty=128; 15'd30922: duty=132; 15'd30923: duty=125; 15'd30924: duty=126; 15'd30925: duty=109; 15'd30926: duty=105; 15'd30927: duty=107;
15'd30928: duty=125; 15'd30929: duty=111; 15'd30930: duty=121; 15'd30931: duty=103; 15'd30932: duty=83; 15'd30933: duty=96; 15'd30934: duty=90; 15'd30935: duty=90;
15'd30936: duty=108; 15'd30937: duty=110; 15'd30938: duty=93; 15'd30939: duty=81; 15'd30940: duty=81; 15'd30941: duty=113; 15'd30942: duty=101; 15'd30943: duty=90;
15'd30944: duty=76; 15'd30945: duty=94; 15'd30946: duty=119; 15'd30947: duty=110; 15'd30948: duty=116; 15'd30949: duty=112; 15'd30950: duty=128; 15'd30951: duty=139;
15'd30952: duty=121; 15'd30953: duty=127; 15'd30954: duty=127; 15'd30955: duty=116; 15'd30956: duty=111; 15'd30957: duty=131; 15'd30958: duty=136; 15'd30959: duty=140;
15'd30960: duty=143; 15'd30961: duty=150; 15'd30962: duty=155; 15'd30963: duty=166; 15'd30964: duty=159; 15'd30965: duty=155; 15'd30966: duty=147; 15'd30967: duty=151;
15'd30968: duty=169; 15'd30969: duty=172; 15'd30970: duty=192; 15'd30971: duty=180; 15'd30972: duty=174; 15'd30973: duty=181; 15'd30974: duty=198; 15'd30975: duty=186;
15'd30976: duty=187; 15'd30977: duty=178; 15'd30978: duty=170; 15'd30979: duty=164; 15'd30980: duty=167; 15'd30981: duty=167; 15'd30982: duty=143; 15'd30983: duty=136;
15'd30984: duty=138; 15'd30985: duty=131; 15'd30986: duty=144; 15'd30987: duty=130; 15'd30988: duty=135; 15'd30989: duty=124; 15'd30990: duty=95; 15'd30991: duty=100;
15'd30992: duty=99; 15'd30993: duty=104; 15'd30994: duty=104; 15'd30995: duty=112; 15'd30996: duty=113; 15'd30997: duty=99; 15'd30998: duty=85; 15'd30999: duty=101;
15'd31000: duty=90; 15'd31001: duty=83; 15'd31002: duty=90; 15'd31003: duty=93; 15'd31004: duty=97; 15'd31005: duty=118; 15'd31006: duty=107; 15'd31007: duty=93;
15'd31008: duty=84; 15'd31009: duty=78; 15'd31010: duty=76; 15'd31011: duty=93; 15'd31012: duty=111; 15'd31013: duty=107; 15'd31014: duty=110; 15'd31015: duty=119;
15'd31016: duty=108; 15'd31017: duty=122; 15'd31018: duty=125; 15'd31019: duty=127; 15'd31020: duty=143; 15'd31021: duty=134; 15'd31022: duty=138; 15'd31023: duty=119;
15'd31024: duty=131; 15'd31025: duty=148; 15'd31026: duty=148; 15'd31027: duty=137; 15'd31028: duty=147; 15'd31029: duty=154; 15'd31030: duty=157; 15'd31031: duty=139;
15'd31032: duty=131; 15'd31033: duty=143; 15'd31034: duty=126; 15'd31035: duty=134; 15'd31036: duty=144; 15'd31037: duty=146; 15'd31038: duty=147; 15'd31039: duty=163;
15'd31040: duty=172; 15'd31041: duty=166; 15'd31042: duty=181; 15'd31043: duty=166; 15'd31044: duty=161; 15'd31045: duty=173; 15'd31046: duty=182; 15'd31047: duty=183;
15'd31048: duty=164; 15'd31049: duty=155; 15'd31050: duty=153; 15'd31051: duty=143; 15'd31052: duty=149; 15'd31053: duty=157; 15'd31054: duty=140; 15'd31055: duty=128;
15'd31056: duty=142; 15'd31057: duty=149; 15'd31058: duty=130; 15'd31059: duty=131; 15'd31060: duty=153; 15'd31061: duty=127; 15'd31062: duty=116; 15'd31063: duty=121;
15'd31064: duty=109; 15'd31065: duty=118; 15'd31066: duty=117; 15'd31067: duty=120; 15'd31068: duty=119; 15'd31069: duty=137; 15'd31070: duty=131; 15'd31071: duty=112;
15'd31072: duty=124; 15'd31073: duty=102; 15'd31074: duty=88; 15'd31075: duty=112; 15'd31076: duty=96; 15'd31077: duty=93; 15'd31078: duty=102; 15'd31079: duty=107;
15'd31080: duty=115; 15'd31081: duty=104; 15'd31082: duty=110; 15'd31083: duty=110; 15'd31084: duty=111; 15'd31085: duty=110; 15'd31086: duty=110; 15'd31087: duty=124;
15'd31088: duty=137; 15'd31089: duty=118; 15'd31090: duty=105; 15'd31091: duty=108; 15'd31092: duty=122; 15'd31093: duty=124; 15'd31094: duty=111; 15'd31095: duty=107;
15'd31096: duty=108; 15'd31097: duty=120; 15'd31098: duty=119; 15'd31099: duty=121; 15'd31100: duty=120; 15'd31101: duty=124; 15'd31102: duty=142; 15'd31103: duty=148;
15'd31104: duty=154; 15'd31105: duty=153; 15'd31106: duty=150; 15'd31107: duty=151; 15'd31108: duty=148; 15'd31109: duty=146; 15'd31110: duty=156; 15'd31111: duty=155;
15'd31112: duty=148; 15'd31113: duty=158; 15'd31114: duty=145; 15'd31115: duty=165; 15'd31116: duty=174; 15'd31117: duty=161; 15'd31118: duty=162; 15'd31119: duty=152;
15'd31120: duty=161; 15'd31121: duty=150; 15'd31122: duty=153; 15'd31123: duty=143; 15'd31124: duty=148; 15'd31125: duty=165; 15'd31126: duty=162; 15'd31127: duty=160;
15'd31128: duty=127; 15'd31129: duty=113; 15'd31130: duty=112; 15'd31131: duty=114; 15'd31132: duty=119; 15'd31133: duty=124; 15'd31134: duty=122; 15'd31135: duty=110;
15'd31136: duty=113; 15'd31137: duty=121; 15'd31138: duty=124; 15'd31139: duty=116; 15'd31140: duty=110; 15'd31141: duty=113; 15'd31142: duty=107; 15'd31143: duty=95;
15'd31144: duty=95; 15'd31145: duty=101; 15'd31146: duty=91; 15'd31147: duty=78; 15'd31148: duty=100; 15'd31149: duty=120; 15'd31150: duty=118; 15'd31151: duty=125;
15'd31152: duty=119; 15'd31153: duty=107; 15'd31154: duty=102; 15'd31155: duty=110; 15'd31156: duty=129; 15'd31157: duty=116; 15'd31158: duty=118; 15'd31159: duty=127;
15'd31160: duty=126; 15'd31161: duty=134; 15'd31162: duty=133; 15'd31163: duty=130; 15'd31164: duty=124; 15'd31165: duty=129; 15'd31166: duty=129; 15'd31167: duty=140;
15'd31168: duty=142; 15'd31169: duty=132; 15'd31170: duty=133; 15'd31171: duty=144; 15'd31172: duty=133; 15'd31173: duty=131; 15'd31174: duty=147; 15'd31175: duty=147;
15'd31176: duty=158; 15'd31177: duty=163; 15'd31178: duty=161; 15'd31179: duty=166; 15'd31180: duty=165; 15'd31181: duty=157; 15'd31182: duty=155; 15'd31183: duty=160;
15'd31184: duty=160; 15'd31185: duty=152; 15'd31186: duty=164; 15'd31187: duty=169; 15'd31188: duty=178; 15'd31189: duty=174; 15'd31190: duty=170; 15'd31191: duty=166;
15'd31192: duty=168; 15'd31193: duty=161; 15'd31194: duty=149; 15'd31195: duty=140; 15'd31196: duty=125; 15'd31197: duty=143; 15'd31198: duty=130; 15'd31199: duty=133;
15'd31200: duty=136; 15'd31201: duty=136; 15'd31202: duty=139; 15'd31203: duty=118; 15'd31204: duty=111; 15'd31205: duty=137; 15'd31206: duty=130; 15'd31207: duty=109;
15'd31208: duty=117; 15'd31209: duty=104; 15'd31210: duty=93; 15'd31211: duty=100; 15'd31212: duty=110; 15'd31213: duty=92; 15'd31214: duty=88; 15'd31215: duty=107;
15'd31216: duty=108; 15'd31217: duty=103; 15'd31218: duty=120; 15'd31219: duty=123; 15'd31220: duty=110; 15'd31221: duty=103; 15'd31222: duty=105; 15'd31223: duty=96;
15'd31224: duty=87; 15'd31225: duty=91; 15'd31226: duty=83; 15'd31227: duty=96; 15'd31228: duty=125; 15'd31229: duty=121; 15'd31230: duty=124; 15'd31231: duty=117;
15'd31232: duty=113; 15'd31233: duty=126; 15'd31234: duty=126; 15'd31235: duty=119; 15'd31236: duty=114; 15'd31237: duty=121; 15'd31238: duty=121; 15'd31239: duty=112;
15'd31240: duty=116; 15'd31241: duty=136; 15'd31242: duty=134; 15'd31243: duty=137; 15'd31244: duty=144; 15'd31245: duty=143; 15'd31246: duty=153; 15'd31247: duty=147;
15'd31248: duty=140; 15'd31249: duty=139; 15'd31250: duty=137; 15'd31251: duty=143; 15'd31252: duty=142; 15'd31253: duty=158; 15'd31254: duty=156; 15'd31255: duty=152;
15'd31256: duty=168; 15'd31257: duty=177; 15'd31258: duty=173; 15'd31259: duty=159; 15'd31260: duty=156; 15'd31261: duty=153; 15'd31262: duty=162; 15'd31263: duty=166;
15'd31264: duty=163; 15'd31265: duty=157; 15'd31266: duty=157; 15'd31267: duty=160; 15'd31268: duty=152; 15'd31269: duty=142; 15'd31270: duty=128; 15'd31271: duty=127;
15'd31272: duty=133; 15'd31273: duty=141; 15'd31274: duty=145; 15'd31275: duty=119; 15'd31276: duty=109; 15'd31277: duty=104; 15'd31278: duty=101; 15'd31279: duty=106;
15'd31280: duty=110; 15'd31281: duty=123; 15'd31282: duty=112; 15'd31283: duty=113; 15'd31284: duty=109; 15'd31285: duty=106; 15'd31286: duty=123; 15'd31287: duty=121;
15'd31288: duty=113; 15'd31289: duty=115; 15'd31290: duty=125; 15'd31291: duty=139; 15'd31292: duty=139; 15'd31293: duty=117; 15'd31294: duty=110; 15'd31295: duty=112;
15'd31296: duty=116; 15'd31297: duty=101; 15'd31298: duty=88; 15'd31299: duty=100; 15'd31300: duty=105; 15'd31301: duty=118; 15'd31302: duty=138; 15'd31303: duty=149;
15'd31304: duty=146; 15'd31305: duty=159; 15'd31306: duty=153; 15'd31307: duty=148; 15'd31308: duty=158; 15'd31309: duty=147; 15'd31310: duty=131; 15'd31311: duty=132;
15'd31312: duty=112; 15'd31313: duty=112; 15'd31314: duty=114; 15'd31315: duty=116; 15'd31316: duty=140; 15'd31317: duty=136; 15'd31318: duty=160; 15'd31319: duty=166;
15'd31320: duty=157; 15'd31321: duty=159; 15'd31322: duty=166; 15'd31323: duty=158; 15'd31324: duty=155; 15'd31325: duty=148; 15'd31326: duty=141; 15'd31327: duty=112;
15'd31328: duty=116; 15'd31329: duty=143; 15'd31330: duty=138; 15'd31331: duty=151; 15'd31332: duty=149; 15'd31333: duty=165; 15'd31334: duty=171; 15'd31335: duty=149;
15'd31336: duty=128; 15'd31337: duty=133; 15'd31338: duty=128; 15'd31339: duty=116; 15'd31340: duty=104; 15'd31341: duty=112; 15'd31342: duty=105; 15'd31343: duty=115;
15'd31344: duty=143; 15'd31345: duty=110; 15'd31346: duty=114; 15'd31347: duty=126; 15'd31348: duty=118; 15'd31349: duty=94; 15'd31350: duty=105; 15'd31351: duty=136;
15'd31352: duty=128; 15'd31353: duty=110; 15'd31354: duty=111; 15'd31355: duty=110; 15'd31356: duty=124; 15'd31357: duty=139; 15'd31358: duty=114; 15'd31359: duty=116;
15'd31360: duty=113; 15'd31361: duty=115; 15'd31362: duty=102; 15'd31363: duty=90; 15'd31364: duty=102; 15'd31365: duty=86; 15'd31366: duty=85; 15'd31367: duty=97;
15'd31368: duty=122; 15'd31369: duty=133; 15'd31370: duty=106; 15'd31371: duty=113; 15'd31372: duty=132; 15'd31373: duty=140; 15'd31374: duty=148; 15'd31375: duty=127;
15'd31376: duty=128; 15'd31377: duty=120; 15'd31378: duty=129; 15'd31379: duty=152; 15'd31380: duty=154; 15'd31381: duty=161; 15'd31382: duty=160; 15'd31383: duty=155;
15'd31384: duty=146; 15'd31385: duty=150; 15'd31386: duty=151; 15'd31387: duty=141; 15'd31388: duty=148; 15'd31389: duty=166; 15'd31390: duty=181; 15'd31391: duty=181;
15'd31392: duty=164; 15'd31393: duty=156; 15'd31394: duty=170; 15'd31395: duty=175; 15'd31396: duty=176; 15'd31397: duty=166; 15'd31398: duty=156; 15'd31399: duty=162;
15'd31400: duty=156; 15'd31401: duty=139; 15'd31402: duty=117; 15'd31403: duty=119; 15'd31404: duty=122; 15'd31405: duty=146; 15'd31406: duty=160; 15'd31407: duty=160;
15'd31408: duty=136; 15'd31409: duty=123; 15'd31410: duty=115; 15'd31411: duty=125; 15'd31412: duty=133; 15'd31413: duty=109; 15'd31414: duty=100; 15'd31415: duty=86;
15'd31416: duty=106; 15'd31417: duty=101; 15'd31418: duty=91; 15'd31419: duty=88; 15'd31420: duty=85; 15'd31421: duty=100; 15'd31422: duty=104; 15'd31423: duty=101;
15'd31424: duty=100; 15'd31425: duty=104; 15'd31426: duty=106; 15'd31427: duty=103; 15'd31428: duty=106; 15'd31429: duty=115; 15'd31430: duty=125; 15'd31431: duty=123;
15'd31432: duty=117; 15'd31433: duty=117; 15'd31434: duty=122; 15'd31435: duty=114; 15'd31436: duty=110; 15'd31437: duty=112; 15'd31438: duty=120; 15'd31439: duty=123;
15'd31440: duty=131; 15'd31441: duty=125; 15'd31442: duty=128; 15'd31443: duty=144; 15'd31444: duty=149; 15'd31445: duty=152; 15'd31446: duty=146; 15'd31447: duty=150;
15'd31448: duty=145; 15'd31449: duty=144; 15'd31450: duty=135; 15'd31451: duty=152; 15'd31452: duty=152; 15'd31453: duty=136; 15'd31454: duty=149; 15'd31455: duty=159;
15'd31456: duty=151; 15'd31457: duty=155; 15'd31458: duty=151; 15'd31459: duty=139; 15'd31460: duty=142; 15'd31461: duty=160; 15'd31462: duty=171; 15'd31463: duty=170;
15'd31464: duty=169; 15'd31465: duty=166; 15'd31466: duty=159; 15'd31467: duty=155; 15'd31468: duty=163; 15'd31469: duty=166; 15'd31470: duty=161; 15'd31471: duty=147;
15'd31472: duty=155; 15'd31473: duty=148; 15'd31474: duty=145; 15'd31475: duty=147; 15'd31476: duty=128; 15'd31477: duty=114; 15'd31478: duty=110; 15'd31479: duty=117;
15'd31480: duty=124; 15'd31481: duty=117; 15'd31482: duty=116; 15'd31483: duty=121; 15'd31484: duty=117; 15'd31485: duty=121; 15'd31486: duty=116; 15'd31487: duty=97;
15'd31488: duty=112; 15'd31489: duty=110; 15'd31490: duty=102; 15'd31491: duty=102; 15'd31492: duty=89; 15'd31493: duty=94; 15'd31494: duty=106; 15'd31495: duty=113;
15'd31496: duty=106; 15'd31497: duty=108; 15'd31498: duty=104; 15'd31499: duty=91; 15'd31500: duty=95; 15'd31501: duty=96; 15'd31502: duty=104; 15'd31503: duty=99;
15'd31504: duty=84; 15'd31505: duty=102; 15'd31506: duty=107; 15'd31507: duty=94; 15'd31508: duty=93; 15'd31509: duty=99; 15'd31510: duty=117; 15'd31511: duty=128;
15'd31512: duty=127; 15'd31513: duty=141; 15'd31514: duty=142; 15'd31515: duty=139; 15'd31516: duty=125; 15'd31517: duty=115; 15'd31518: duty=141; 15'd31519: duty=145;
15'd31520: duty=142; 15'd31521: duty=133; 15'd31522: duty=130; 15'd31523: duty=141; 15'd31524: duty=153; 15'd31525: duty=165; 15'd31526: duty=157; 15'd31527: duty=153;
15'd31528: duty=154; 15'd31529: duty=156; 15'd31530: duty=163; 15'd31531: duty=162; 15'd31532: duty=160; 15'd31533: duty=163; 15'd31534: duty=164; 15'd31535: duty=173;
15'd31536: duty=174; 15'd31537: duty=169; 15'd31538: duty=171; 15'd31539: duty=165; 15'd31540: duty=159; 15'd31541: duty=171; 15'd31542: duty=183; 15'd31543: duty=167;
15'd31544: duty=143; 15'd31545: duty=145; 15'd31546: duty=154; 15'd31547: duty=149; 15'd31548: duty=154; 15'd31549: duty=162; 15'd31550: duty=134; 15'd31551: duty=127;
15'd31552: duty=128; 15'd31553: duty=117; 15'd31554: duty=114; 15'd31555: duty=112; 15'd31556: duty=104; 15'd31557: duty=103; 15'd31558: duty=117; 15'd31559: duty=124;
15'd31560: duty=125; 15'd31561: duty=118; 15'd31562: duty=116; 15'd31563: duty=112; 15'd31564: duty=113; 15'd31565: duty=121; 15'd31566: duty=114; 15'd31567: duty=99;
15'd31568: duty=102; 15'd31569: duty=107; 15'd31570: duty=99; 15'd31571: duty=89; 15'd31572: duty=106; 15'd31573: duty=116; 15'd31574: duty=102; 15'd31575: duty=99;
15'd31576: duty=103; 15'd31577: duty=106; 15'd31578: duty=107; 15'd31579: duty=109; 15'd31580: duty=105; 15'd31581: duty=119; 15'd31582: duty=129; 15'd31583: duty=139;
15'd31584: duty=131; 15'd31585: duty=136; 15'd31586: duty=135; 15'd31587: duty=127; 15'd31588: duty=127; 15'd31589: duty=130; 15'd31590: duty=148; 15'd31591: duty=145;
15'd31592: duty=124; 15'd31593: duty=121; 15'd31594: duty=117; 15'd31595: duty=112; 15'd31596: duty=132; 15'd31597: duty=128; 15'd31598: duty=134; 15'd31599: duty=137;
15'd31600: duty=145; 15'd31601: duty=150; 15'd31602: duty=157; 15'd31603: duty=164; 15'd31604: duty=157; 15'd31605: duty=170; 15'd31606: duty=159; 15'd31607: duty=144;
15'd31608: duty=146; 15'd31609: duty=153; 15'd31610: duty=157; 15'd31611: duty=145; 15'd31612: duty=143; 15'd31613: duty=147; 15'd31614: duty=158; 15'd31615: duty=172;
15'd31616: duty=155; 15'd31617: duty=131; 15'd31618: duty=113; 15'd31619: duty=114; 15'd31620: duty=126; 15'd31621: duty=131; 15'd31622: duty=135; 15'd31623: duty=129;
15'd31624: duty=113; 15'd31625: duty=107; 15'd31626: duty=104; 15'd31627: duty=116; 15'd31628: duty=120; 15'd31629: duty=120; 15'd31630: duty=130; 15'd31631: duty=117;
15'd31632: duty=123; 15'd31633: duty=138; 15'd31634: duty=123; 15'd31635: duty=111; 15'd31636: duty=118; 15'd31637: duty=114; 15'd31638: duty=115; 15'd31639: duty=111;
15'd31640: duty=108; 15'd31641: duty=101; 15'd31642: duty=100; 15'd31643: duty=110; 15'd31644: duty=101; 15'd31645: duty=103; 15'd31646: duty=115; 15'd31647: duty=130;
15'd31648: duty=118; 15'd31649: duty=122; 15'd31650: duty=141; 15'd31651: duty=147; 15'd31652: duty=133; 15'd31653: duty=120; 15'd31654: duty=126; 15'd31655: duty=126;
15'd31656: duty=126; 15'd31657: duty=139; 15'd31658: duty=148; 15'd31659: duty=138; 15'd31660: duty=151; 15'd31661: duty=151; 15'd31662: duty=138; 15'd31663: duty=146;
15'd31664: duty=155; 15'd31665: duty=147; 15'd31666: duty=153; 15'd31667: duty=157; 15'd31668: duty=156; 15'd31669: duty=162; 15'd31670: duty=156; 15'd31671: duty=142;
15'd31672: duty=156; 15'd31673: duty=163; 15'd31674: duty=154; 15'd31675: duty=154; 15'd31676: duty=156; 15'd31677: duty=157; 15'd31678: duty=147; 15'd31679: duty=151;
15'd31680: duty=156; 15'd31681: duty=152; 15'd31682: duty=135; 15'd31683: duty=129; 15'd31684: duty=133; 15'd31685: duty=140; 15'd31686: duty=148; 15'd31687: duty=139;
15'd31688: duty=130; 15'd31689: duty=131; 15'd31690: duty=137; 15'd31691: duty=131; 15'd31692: duty=126; 15'd31693: duty=122; 15'd31694: duty=107; 15'd31695: duty=95;
15'd31696: duty=95; 15'd31697: duty=92; 15'd31698: duty=99; 15'd31699: duty=96; 15'd31700: duty=96; 15'd31701: duty=112; 15'd31702: duty=110; 15'd31703: duty=112;
15'd31704: duty=107; 15'd31705: duty=110; 15'd31706: duty=110; 15'd31707: duty=103; 15'd31708: duty=96; 15'd31709: duty=95; 15'd31710: duty=100; 15'd31711: duty=96;
15'd31712: duty=102; 15'd31713: duty=113; 15'd31714: duty=100; 15'd31715: duty=98; 15'd31716: duty=104; 15'd31717: duty=100; 15'd31718: duty=107; 15'd31719: duty=101;
15'd31720: duty=104; 15'd31721: duty=109; 15'd31722: duty=118; 15'd31723: duty=128; 15'd31724: duty=142; 15'd31725: duty=144; 15'd31726: duty=142; 15'd31727: duty=137;
15'd31728: duty=131; 15'd31729: duty=139; 15'd31730: duty=146; 15'd31731: duty=142; 15'd31732: duty=147; 15'd31733: duty=142; 15'd31734: duty=154; 15'd31735: duty=159;
15'd31736: duty=154; 15'd31737: duty=159; 15'd31738: duty=163; 15'd31739: duty=161; 15'd31740: duty=171; 15'd31741: duty=182; 15'd31742: duty=175; 15'd31743: duty=173;
15'd31744: duty=178; 15'd31745: duty=187; 15'd31746: duty=168; 15'd31747: duty=176; 15'd31748: duty=163; 15'd31749: duty=159; 15'd31750: duty=163; 15'd31751: duty=162;
15'd31752: duty=166; 15'd31753: duty=162; 15'd31754: duty=155; 15'd31755: duty=164; 15'd31756: duty=162; 15'd31757: duty=148; 15'd31758: duty=140; 15'd31759: duty=142;
15'd31760: duty=134; 15'd31761: duty=120; 15'd31762: duty=134; 15'd31763: duty=128; 15'd31764: duty=136; 15'd31765: duty=127; 15'd31766: duty=120; 15'd31767: duty=107;
15'd31768: duty=90; 15'd31769: duty=99; 15'd31770: duty=91; 15'd31771: duty=93; 15'd31772: duty=89; 15'd31773: duty=88; 15'd31774: duty=115; 15'd31775: duty=110;
15'd31776: duty=110; 15'd31777: duty=91; 15'd31778: duty=81; 15'd31779: duty=87; 15'd31780: duty=95; 15'd31781: duty=109; 15'd31782: duty=99; 15'd31783: duty=98;
15'd31784: duty=98; 15'd31785: duty=91; 15'd31786: duty=95; 15'd31787: duty=88; 15'd31788: duty=94; 15'd31789: duty=96; 15'd31790: duty=107; 15'd31791: duty=124;
15'd31792: duty=124; 15'd31793: duty=137; 15'd31794: duty=123; 15'd31795: duty=129; 15'd31796: duty=115; 15'd31797: duty=128; 15'd31798: duty=149; 15'd31799: duty=140;
15'd31800: duty=139; 15'd31801: duty=140; 15'd31802: duty=147; 15'd31803: duty=151; 15'd31804: duty=142; 15'd31805: duty=132; 15'd31806: duty=147; 15'd31807: duty=168;
15'd31808: duty=172; 15'd31809: duty=147; 15'd31810: duty=141; 15'd31811: duty=165; 15'd31812: duty=163; 15'd31813: duty=146; 15'd31814: duty=151; 15'd31815: duty=171;
15'd31816: duty=173; 15'd31817: duty=156; 15'd31818: duty=160; 15'd31819: duty=165; 15'd31820: duty=160; 15'd31821: duty=161; 15'd31822: duty=159; 15'd31823: duty=159;
15'd31824: duty=165; 15'd31825: duty=159; 15'd31826: duty=154; 15'd31827: duty=138; 15'd31828: duty=128; 15'd31829: duty=130; 15'd31830: duty=131; 15'd31831: duty=121;
15'd31832: duty=131; 15'd31833: duty=138; 15'd31834: duty=117; 15'd31835: duty=126; 15'd31836: duty=125; 15'd31837: duty=119; 15'd31838: duty=119; 15'd31839: duty=107;
15'd31840: duty=107; 15'd31841: duty=107; 15'd31842: duty=96; 15'd31843: duty=97; 15'd31844: duty=103; 15'd31845: duty=99; 15'd31846: duty=93; 15'd31847: duty=98;
15'd31848: duty=94; 15'd31849: duty=101; 15'd31850: duty=111; 15'd31851: duty=107; 15'd31852: duty=105; 15'd31853: duty=109; 15'd31854: duty=108; 15'd31855: duty=100;
15'd31856: duty=99; 15'd31857: duty=103; 15'd31858: duty=107; 15'd31859: duty=106; 15'd31860: duty=110; 15'd31861: duty=99; 15'd31862: duty=102; 15'd31863: duty=127;
15'd31864: duty=143; 15'd31865: duty=142; 15'd31866: duty=149; 15'd31867: duty=136; 15'd31868: duty=131; 15'd31869: duty=148; 15'd31870: duty=147; 15'd31871: duty=149;
15'd31872: duty=138; 15'd31873: duty=136; 15'd31874: duty=123; 15'd31875: duty=130; 15'd31876: duty=160; 15'd31877: duty=142; 15'd31878: duty=129; 15'd31879: duty=136;
15'd31880: duty=151; 15'd31881: duty=167; 15'd31882: duty=171; 15'd31883: duty=163; 15'd31884: duty=169; 15'd31885: duty=190; 15'd31886: duty=184; 15'd31887: duty=176;
15'd31888: duty=162; 15'd31889: duty=152; 15'd31890: duty=168; 15'd31891: duty=165; 15'd31892: duty=157; 15'd31893: duty=174; 15'd31894: duty=182; 15'd31895: duty=176;
15'd31896: duty=153; 15'd31897: duty=143; 15'd31898: duty=162; 15'd31899: duty=144; 15'd31900: duty=133; 15'd31901: duty=132; 15'd31902: duty=122; 15'd31903: duty=145;
15'd31904: duty=141; 15'd31905: duty=130; 15'd31906: duty=126; 15'd31907: duty=125; 15'd31908: duty=128; 15'd31909: duty=116; 15'd31910: duty=132; 15'd31911: duty=121;
15'd31912: duty=101; 15'd31913: duty=110; 15'd31914: duty=93; 15'd31915: duty=97; 15'd31916: duty=104; 15'd31917: duty=89; 15'd31918: duty=90; 15'd31919: duty=85;
15'd31920: duty=84; 15'd31921: duty=86; 15'd31922: duty=107; 15'd31923: duty=118; 15'd31924: duty=107; 15'd31925: duty=101; 15'd31926: duty=86; 15'd31927: duty=90;
15'd31928: duty=98; 15'd31929: duty=102; 15'd31930: duty=84; 15'd31931: duty=89; 15'd31932: duty=116; 15'd31933: duty=118; 15'd31934: duty=102; 15'd31935: duty=102;
15'd31936: duty=108; 15'd31937: duty=104; 15'd31938: duty=111; 15'd31939: duty=104; 15'd31940: duty=123; 15'd31941: duty=139; 15'd31942: duty=125; 15'd31943: duty=118;
15'd31944: duty=136; 15'd31945: duty=155; 15'd31946: duty=161; 15'd31947: duty=154; 15'd31948: duty=138; 15'd31949: duty=151; 15'd31950: duty=169; 15'd31951: duty=154;
15'd31952: duty=150; 15'd31953: duty=150; 15'd31954: duty=158; 15'd31955: duty=166; 15'd31956: duty=168; 15'd31957: duty=173; 15'd31958: duty=160; 15'd31959: duty=162;
15'd31960: duty=171; 15'd31961: duty=153; 15'd31962: duty=171; 15'd31963: duty=181; 15'd31964: duty=163; 15'd31965: duty=157; 15'd31966: duty=157; 15'd31967: duty=170;
15'd31968: duty=171; 15'd31969: duty=153; 15'd31970: duty=142; 15'd31971: duty=145; 15'd31972: duty=145; 15'd31973: duty=142; 15'd31974: duty=128; 15'd31975: duty=133;
15'd31976: duty=112; 15'd31977: duty=107; 15'd31978: duty=111; 15'd31979: duty=119; 15'd31980: duty=121; 15'd31981: duty=96; 15'd31982: duty=110; 15'd31983: duty=102;
15'd31984: duty=95; 15'd31985: duty=125; 15'd31986: duty=109; 15'd31987: duty=100; 15'd31988: duty=101; 15'd31989: duty=95; 15'd31990: duty=110; 15'd31991: duty=95;
15'd31992: duty=106; 15'd31993: duty=110; 15'd31994: duty=115; 15'd31995: duty=114; 15'd31996: duty=90; 15'd31997: duty=88; 15'd31998: duty=91; 15'd31999: duty=89;
15'd32000: duty=115; 15'd32001: duty=128; 15'd32002: duty=134; 15'd32003: duty=146; 15'd32004: duty=150; 15'd32005: duty=155; 15'd32006: duty=156; 15'd32007: duty=143;
15'd32008: duty=126; 15'd32009: duty=122; 15'd32010: duty=124; 15'd32011: duty=142; 15'd32012: duty=150; 15'd32013: duty=151; 15'd32014: duty=124; 15'd32015: duty=135;
15'd32016: duty=146; 15'd32017: duty=143; 15'd32018: duty=145; 15'd32019: duty=153; 15'd32020: duty=143; 15'd32021: duty=139; 15'd32022: duty=145; 15'd32023: duty=148;
15'd32024: duty=143; 15'd32025: duty=150; 15'd32026: duty=165; 15'd32027: duty=150; 15'd32028: duty=153; 15'd32029: duty=167; 15'd32030: duty=171; 15'd32031: duty=164;
15'd32032: duty=163; 15'd32033: duty=159; 15'd32034: duty=167; 15'd32035: duty=161; 15'd32036: duty=152; 15'd32037: duty=130; 15'd32038: duty=126; 15'd32039: duty=134;
15'd32040: duty=131; 15'd32041: duty=111; 15'd32042: duty=126; 15'd32043: duty=138; 15'd32044: duty=117; 15'd32045: duty=106; 15'd32046: duty=127; 15'd32047: duty=126;
15'd32048: duty=108; 15'd32049: duty=102; 15'd32050: duty=94; 15'd32051: duty=123; 15'd32052: duty=117; 15'd32053: duty=96; 15'd32054: duty=106; 15'd32055: duty=121;
15'd32056: duty=116; 15'd32057: duty=114; 15'd32058: duty=99; 15'd32059: duty=107; 15'd32060: duty=116; 15'd32061: duty=115; 15'd32062: duty=103; 15'd32063: duty=88;
15'd32064: duty=101; 15'd32065: duty=87; 15'd32066: duty=80; 15'd32067: duty=106; 15'd32068: duty=109; 15'd32069: duty=92; 15'd32070: duty=89; 15'd32071: duty=104;
15'd32072: duty=119; 15'd32073: duty=121; 15'd32074: duty=143; 15'd32075: duty=133; 15'd32076: duty=116; 15'd32077: duty=126; 15'd32078: duty=129; 15'd32079: duty=124;
15'd32080: duty=114; 15'd32081: duty=130; 15'd32082: duty=126; 15'd32083: duty=142; 15'd32084: duty=139; 15'd32085: duty=130; 15'd32086: duty=157; 15'd32087: duty=161;
15'd32088: duty=159; 15'd32089: duty=158; 15'd32090: duty=143; 15'd32091: duty=148; 15'd32092: duty=168; 15'd32093: duty=161; 15'd32094: duty=166; 15'd32095: duty=171;
15'd32096: duty=197; 15'd32097: duty=180; 15'd32098: duty=162; 15'd32099: duty=168; 15'd32100: duty=173; 15'd32101: duty=182; 15'd32102: duty=180; 15'd32103: duty=159;
15'd32104: duty=182; 15'd32105: duty=193; 15'd32106: duty=175; 15'd32107: duty=171; 15'd32108: duty=156; 15'd32109: duty=153; 15'd32110: duty=139; 15'd32111: duty=128;
15'd32112: duty=121; 15'd32113: duty=140; 15'd32114: duty=140; 15'd32115: duty=128; 15'd32116: duty=128; 15'd32117: duty=109; 15'd32118: duty=118; 15'd32119: duty=128;
15'd32120: duty=95; 15'd32121: duty=95; 15'd32122: duty=107; 15'd32123: duty=113; 15'd32124: duty=118; 15'd32125: duty=105; 15'd32126: duty=117; 15'd32127: duty=135;
15'd32128: duty=109; 15'd32129: duty=96; 15'd32130: duty=83; 15'd32131: duty=87; 15'd32132: duty=91; 15'd32133: duty=95; 15'd32134: duty=108; 15'd32135: duty=99;
15'd32136: duty=105; 15'd32137: duty=92; 15'd32138: duty=100; 15'd32139: duty=98; 15'd32140: duty=94; 15'd32141: duty=106; 15'd32142: duty=93; 15'd32143: duty=119;
15'd32144: duty=129; 15'd32145: duty=96; 15'd32146: duty=122; 15'd32147: duty=146; 15'd32148: duty=130; 15'd32149: duty=123; 15'd32150: duty=127; 15'd32151: duty=129;
15'd32152: duty=125; 15'd32153: duty=129; 15'd32154: duty=125; 15'd32155: duty=117; 15'd32156: duty=127; 15'd32157: duty=119; 15'd32158: duty=123; 15'd32159: duty=128;
15'd32160: duty=123; 15'd32161: duty=145; 15'd32162: duty=137; 15'd32163: duty=134; 15'd32164: duty=145; 15'd32165: duty=146; 15'd32166: duty=154; 15'd32167: duty=155;
15'd32168: duty=132; 15'd32169: duty=127; 15'd32170: duty=152; 15'd32171: duty=158; 15'd32172: duty=171; 15'd32173: duty=170; 15'd32174: duty=162; 15'd32175: duty=160;
15'd32176: duty=156; 15'd32177: duty=161; 15'd32178: duty=160; 15'd32179: duty=148; 15'd32180: duty=137; 15'd32181: duty=127; 15'd32182: duty=119; 15'd32183: duty=122;
15'd32184: duty=135; 15'd32185: duty=150; 15'd32186: duty=141; 15'd32187: duty=133; 15'd32188: duty=147; 15'd32189: duty=157; 15'd32190: duty=154; 15'd32191: duty=135;
15'd32192: duty=116; 15'd32193: duty=118; 15'd32194: duty=120; 15'd32195: duty=131; 15'd32196: duty=138; 15'd32197: duty=131; 15'd32198: duty=123; 15'd32199: duty=121;
15'd32200: duty=123; 15'd32201: duty=138; 15'd32202: duty=152; 15'd32203: duty=139; 15'd32204: duty=121; 15'd32205: duty=132; 15'd32206: duty=138; 15'd32207: duty=126;
15'd32208: duty=117; 15'd32209: duty=108; 15'd32210: duty=118; 15'd32211: duty=120; 15'd32212: duty=108; 15'd32213: duty=103; 15'd32214: duty=118; 15'd32215: duty=134;
15'd32216: duty=144; 15'd32217: duty=119; 15'd32218: duty=117; 15'd32219: duty=128; 15'd32220: duty=126; 15'd32221: duty=126; 15'd32222: duty=110; 15'd32223: duty=129;
15'd32224: duty=142; 15'd32225: duty=131; 15'd32226: duty=129; 15'd32227: duty=137; 15'd32228: duty=135; 15'd32229: duty=129; 15'd32230: duty=128; 15'd32231: duty=131;
15'd32232: duty=127; 15'd32233: duty=130; 15'd32234: duty=141; 15'd32235: duty=131; 15'd32236: duty=130; 15'd32237: duty=137; 15'd32238: duty=146; 15'd32239: duty=143;
15'd32240: duty=136; 15'd32241: duty=146; 15'd32242: duty=145; 15'd32243: duty=145; 15'd32244: duty=142; 15'd32245: duty=142; 15'd32246: duty=145; 15'd32247: duty=134;
15'd32248: duty=131; 15'd32249: duty=118; 15'd32250: duty=132; 15'd32251: duty=137; 15'd32252: duty=136; 15'd32253: duty=122; 15'd32254: duty=115; 15'd32255: duty=122;
15'd32256: duty=115; 15'd32257: duty=112; 15'd32258: duty=105; 15'd32259: duty=125; 15'd32260: duty=107; 15'd32261: duty=119; 15'd32262: duty=110; 15'd32263: duty=99;
15'd32264: duty=115; 15'd32265: duty=110; 15'd32266: duty=120; 15'd32267: duty=119; 15'd32268: duty=123; 15'd32269: duty=113; 15'd32270: duty=118; 15'd32271: duty=122;
15'd32272: duty=115; 15'd32273: duty=119; 15'd32274: duty=106; 15'd32275: duty=111; 15'd32276: duty=112; 15'd32277: duty=97; 15'd32278: duty=106; 15'd32279: duty=115;
15'd32280: duty=121; 15'd32281: duty=131; 15'd32282: duty=139; 15'd32283: duty=160; 15'd32284: duty=156; 15'd32285: duty=140; 15'd32286: duty=140; 15'd32287: duty=157;
15'd32288: duty=156; 15'd32289: duty=139; 15'd32290: duty=128; 15'd32291: duty=121; 15'd32292: duty=140; 15'd32293: duty=150; 15'd32294: duty=150; 15'd32295: duty=121;
15'd32296: duty=141; 15'd32297: duty=151; 15'd32298: duty=151; 15'd32299: duty=145; 15'd32300: duty=144; 15'd32301: duty=160; 15'd32302: duty=144; 15'd32303: duty=145;
15'd32304: duty=154; 15'd32305: duty=174; 15'd32306: duty=171; 15'd32307: duty=163; 15'd32308: duty=147; 15'd32309: duty=155; 15'd32310: duty=165; 15'd32311: duty=158;
15'd32312: duty=152; 15'd32313: duty=164; 15'd32314: duty=170; 15'd32315: duty=169; 15'd32316: duty=160; 15'd32317: duty=149; 15'd32318: duty=162; 15'd32319: duty=155;
15'd32320: duty=139; 15'd32321: duty=134; 15'd32322: duty=135; 15'd32323: duty=141; 15'd32324: duty=136; 15'd32325: duty=102; 15'd32326: duty=102; 15'd32327: duty=115;
15'd32328: duty=136; 15'd32329: duty=146; 15'd32330: duty=124; 15'd32331: duty=113; 15'd32332: duty=112; 15'd32333: duty=125; 15'd32334: duty=106; 15'd32335: duty=95;
15'd32336: duty=92; 15'd32337: duty=90; 15'd32338: duty=80; 15'd32339: duty=93; 15'd32340: duty=116; 15'd32341: duty=116; 15'd32342: duty=107; 15'd32343: duty=101;
15'd32344: duty=101; 15'd32345: duty=95; 15'd32346: duty=93; 15'd32347: duty=82; 15'd32348: duty=79; 15'd32349: duty=61; 15'd32350: duty=75; 15'd32351: duty=97;
15'd32352: duty=82; 15'd32353: duty=92; 15'd32354: duty=115; 15'd32355: duty=114; 15'd32356: duty=111; 15'd32357: duty=112; 15'd32358: duty=105; 15'd32359: duty=110;
15'd32360: duty=113; 15'd32361: duty=110; 15'd32362: duty=121; 15'd32363: duty=133; 15'd32364: duty=156; 15'd32365: duty=154; 15'd32366: duty=145; 15'd32367: duty=161;
15'd32368: duty=156; 15'd32369: duty=151; 15'd32370: duty=168; 15'd32371: duty=153; 15'd32372: duty=157; 15'd32373: duty=158; 15'd32374: duty=157; 15'd32375: duty=168;
15'd32376: duty=157; 15'd32377: duty=170; 15'd32378: duty=165; 15'd32379: duty=164; 15'd32380: duty=171; 15'd32381: duty=185; 15'd32382: duty=197; 15'd32383: duty=201;
15'd32384: duty=191; 15'd32385: duty=171; 15'd32386: duty=149; 15'd32387: duty=148; 15'd32388: duty=148; 15'd32389: duty=137; 15'd32390: duty=143; 15'd32391: duty=132;
15'd32392: duty=134; 15'd32393: duty=155; 15'd32394: duty=132; 15'd32395: duty=123; 15'd32396: duty=115; 15'd32397: duty=128; 15'd32398: duty=145; 15'd32399: duty=129;
15'd32400: duty=126; 15'd32401: duty=121; 15'd32402: duty=108; 15'd32403: duty=104; 15'd32404: duty=124; 15'd32405: duty=121; 15'd32406: duty=122; 15'd32407: duty=116;
15'd32408: duty=95; 15'd32409: duty=96; 15'd32410: duty=109; 15'd32411: duty=120; 15'd32412: duty=104; 15'd32413: duty=89; 15'd32414: duty=108; 15'd32415: duty=114;
15'd32416: duty=125; 15'd32417: duty=124; 15'd32418: duty=123; 15'd32419: duty=113; 15'd32420: duty=95; 15'd32421: duty=112; 15'd32422: duty=120; 15'd32423: duty=111;
15'd32424: duty=110; 15'd32425: duty=108; 15'd32426: duty=124; 15'd32427: duty=128; 15'd32428: duty=136; 15'd32429: duty=152; 15'd32430: duty=114; 15'd32431: duty=121;
15'd32432: duty=137; 15'd32433: duty=134; 15'd32434: duty=142; 15'd32435: duty=134; 15'd32436: duty=123; 15'd32437: duty=121; 15'd32438: duty=130; 15'd32439: duty=139;
15'd32440: duty=128; 15'd32441: duty=131; 15'd32442: duty=127; 15'd32443: duty=128; 15'd32444: duty=147; 15'd32445: duty=157; 15'd32446: duty=152; 15'd32447: duty=140;
15'd32448: duty=134; 15'd32449: duty=139; 15'd32450: duty=169; 15'd32451: duty=166; 15'd32452: duty=143; 15'd32453: duty=128; 15'd32454: duty=130; 15'd32455: duty=143;
15'd32456: duty=164; 15'd32457: duty=153; 15'd32458: duty=139; 15'd32459: duty=142; 15'd32460: duty=139; 15'd32461: duty=133; 15'd32462: duty=129; 15'd32463: duty=137;
15'd32464: duty=119; 15'd32465: duty=110; 15'd32466: duty=134; 15'd32467: duty=139; 15'd32468: duty=134; 15'd32469: duty=140; 15'd32470: duty=118; 15'd32471: duty=128;
15'd32472: duty=131; 15'd32473: duty=118; 15'd32474: duty=131; 15'd32475: duty=124; 15'd32476: duty=130; 15'd32477: duty=125; 15'd32478: duty=111; 15'd32479: duty=118;
15'd32480: duty=105; 15'd32481: duty=117; 15'd32482: duty=118; 15'd32483: duty=104; 15'd32484: duty=111; 15'd32485: duty=115; 15'd32486: duty=132; 15'd32487: duty=134;
15'd32488: duty=124; 15'd32489: duty=111; 15'd32490: duty=108; 15'd32491: duty=116; 15'd32492: duty=124; 15'd32493: duty=118; 15'd32494: duty=114; 15'd32495: duty=114;
15'd32496: duty=123; 15'd32497: duty=124; 15'd32498: duty=114; 15'd32499: duty=126; 15'd32500: duty=127; 15'd32501: duty=130; 15'd32502: duty=131; 15'd32503: duty=133;
15'd32504: duty=145; 15'd32505: duty=147; 15'd32506: duty=145; 15'd32507: duty=161; 15'd32508: duty=168; 15'd32509: duty=154; 15'd32510: duty=153; 15'd32511: duty=161;
15'd32512: duty=157; 15'd32513: duty=155; 15'd32514: duty=163; 15'd32515: duty=159; 15'd32516: duty=146; 15'd32517: duty=138; 15'd32518: duty=149; 15'd32519: duty=165;
15'd32520: duty=154; 15'd32521: duty=154; 15'd32522: duty=160; 15'd32523: duty=162; 15'd32524: duty=153; 15'd32525: duty=134; 15'd32526: duty=142; 15'd32527: duty=139;
15'd32528: duty=121; 15'd32529: duty=141; 15'd32530: duty=139; 15'd32531: duty=115; 15'd32532: duty=111; 15'd32533: duty=114; 15'd32534: duty=127; 15'd32535: duty=104;
15'd32536: duty=107; 15'd32537: duty=104; 15'd32538: duty=91; 15'd32539: duty=95; 15'd32540: duty=101; 15'd32541: duty=113; 15'd32542: duty=105; 15'd32543: duty=98;
15'd32544: duty=94; 15'd32545: duty=105; 15'd32546: duty=96; 15'd32547: duty=94; 15'd32548: duty=99; 15'd32549: duty=101; 15'd32550: duty=93; 15'd32551: duty=87;
15'd32552: duty=96; 15'd32553: duty=102; 15'd32554: duty=113; 15'd32555: duty=113; 15'd32556: duty=96; 15'd32557: duty=93; 15'd32558: duty=110; 15'd32559: duty=132;
15'd32560: duty=134; 15'd32561: duty=145; 15'd32562: duty=156; 15'd32563: duty=147; 15'd32564: duty=148; 15'd32565: duty=149; 15'd32566: duty=169; 15'd32567: duty=171;
15'd32568: duty=162; 15'd32569: duty=162; 15'd32570: duty=154; 15'd32571: duty=149; 15'd32572: duty=158; 15'd32573: duty=154; 15'd32574: duty=145; 15'd32575: duty=137;
15'd32576: duty=131; 15'd32577: duty=151; 15'd32578: duty=162; 15'd32579: duty=161; 15'd32580: duty=167; 15'd32581: duty=157; 15'd32582: duty=149; 15'd32583: duty=160;
15'd32584: duty=158; 15'd32585: duty=157; 15'd32586: duty=167; 15'd32587: duty=152; 15'd32588: duty=147; 15'd32589: duty=149; 15'd32590: duty=147; 15'd32591: duty=155;
15'd32592: duty=160; 15'd32593: duty=159; 15'd32594: duty=151; 15'd32595: duty=154; 15'd32596: duty=159; 15'd32597: duty=146; 15'd32598: duty=130; 15'd32599: duty=134;
15'd32600: duty=109; 15'd32601: duty=104; 15'd32602: duty=101; 15'd32603: duty=96; 15'd32604: duty=116; 15'd32605: duty=105; 15'd32606: duty=93; 15'd32607: duty=101;
15'd32608: duty=109; 15'd32609: duty=106; 15'd32610: duty=99; 15'd32611: duty=95; 15'd32612: duty=107; 15'd32613: duty=101; 15'd32614: duty=81; 15'd32615: duty=90;
15'd32616: duty=102; 15'd32617: duty=106; 15'd32618: duty=107; 15'd32619: duty=103; 15'd32620: duty=109; 15'd32621: duty=109; 15'd32622: duty=112; 15'd32623: duty=126;
15'd32624: duty=120; 15'd32625: duty=86; 15'd32626: duty=87; 15'd32627: duty=100; 15'd32628: duty=100; 15'd32629: duty=123; 15'd32630: duty=121; 15'd32631: duty=115;
15'd32632: duty=125; 15'd32633: duty=144; 15'd32634: duty=153; 15'd32635: duty=156; 15'd32636: duty=144; 15'd32637: duty=131; 15'd32638: duty=135; 15'd32639: duty=153;
15'd32640: duty=168; 15'd32641: duty=160; 15'd32642: duty=151; 15'd32643: duty=137; 15'd32644: duty=134; 15'd32645: duty=151; 15'd32646: duty=168; 15'd32647: duty=176;
15'd32648: duty=166; 15'd32649: duty=151; 15'd32650: duty=162; 15'd32651: duty=165; 15'd32652: duty=153; 15'd32653: duty=139; 15'd32654: duty=159; 15'd32655: duty=164;
15'd32656: duty=154; 15'd32657: duty=162; 15'd32658: duty=164; 15'd32659: duty=174; 15'd32660: duty=179; 15'd32661: duty=165; 15'd32662: duty=154; 15'd32663: duty=157;
15'd32664: duty=162; 15'd32665: duty=154; 15'd32666: duty=121; 15'd32667: duty=141; 15'd32668: duty=156; 15'd32669: duty=127; 15'd32670: duty=107; 15'd32671: duty=117;
15'd32672: duty=123; 15'd32673: duty=122; 15'd32674: duty=104; 15'd32675: duty=100; 15'd32676: duty=119; 15'd32677: duty=99; 15'd32678: duty=102; 15'd32679: duty=95;
15'd32680: duty=107; 15'd32681: duty=105; 15'd32682: duty=85; 15'd32683: duty=84; 15'd32684: duty=87; 15'd32685: duty=97; 15'd32686: duty=92; 15'd32687: duty=71;
15'd32688: duty=79; 15'd32689: duty=95; 15'd32690: duty=104; 15'd32691: duty=113; 15'd32692: duty=99; 15'd32693: duty=100; 15'd32694: duty=99; 15'd32695: duty=106;
15'd32696: duty=122; 15'd32697: duty=113; 15'd32698: duty=111; 15'd32699: duty=116; 15'd32700: duty=115; 15'd32701: duty=123; 15'd32702: duty=122; 15'd32703: duty=134;
15'd32704: duty=136; 15'd32705: duty=137; 15'd32706: duty=144; 15'd32707: duty=149; 15'd32708: duty=150; 15'd32709: duty=134; 15'd32710: duty=137; 15'd32711: duty=154;
15'd32712: duty=156; 15'd32713: duty=160; 15'd32714: duty=171; 15'd32715: duty=166; 15'd32716: duty=153; 15'd32717: duty=149; 15'd32718: duty=146; 15'd32719: duty=143;
15'd32720: duty=162; 15'd32721: duty=157; 15'd32722: duty=160; 15'd32723: duty=174; 15'd32724: duty=171; 15'd32725: duty=160; 15'd32726: duty=162; 15'd32727: duty=173;
15'd32728: duty=157; 15'd32729: duty=154; 15'd32730: duty=158; 15'd32731: duty=159; 15'd32732: duty=154; 15'd32733: duty=157; 15'd32734: duty=160; 15'd32735: duty=146;
15'd32736: duty=132; 15'd32737: duty=121; 15'd32738: duty=149; 15'd32739: duty=132; 15'd32740: duty=114; 15'd32741: duty=129; 15'd32742: duty=117; 15'd32743: duty=113;
15'd32744: duty=114; 15'd32745: duty=120; 15'd32746: duty=113; 15'd32747: duty=115; 15'd32748: duty=131; 15'd32749: duty=114; 15'd32750: duty=93; 15'd32751: duty=106;
15'd32752: duty=126; 15'd32753: duty=130; 15'd32754: duty=91; 15'd32755: duty=83; 15'd32756: duty=97; 15'd32757: duty=81; 15'd32758: duty=74; 15'd32759: duty=80;
15'd32760: duty=100; 15'd32761: duty=107; 15'd32762: duty=97; 15'd32763: duty=81; 15'd32764: duty=105; 15'd32765: duty=118; 15'd32766: duty=121; 15'd32767: duty=124;



default: duty = 0;
endcase


endmodule
